library ieee;
use ieee.std_logic_1164.all;
use work.my_package.all;
-----------------------------------------------
entity CUTs is
	generic(
		g_N_Segments	:	integer;
		g_N_Parallel	:	integer
	);
	port(
		i_Clk_Launch	:	in	std_logic;
		i_Clk_Sample	:	in	std_logic;
		i_CE	:	in	std_logic;
		i_CLR	:	in	std_logic;
		o_Error	:	out	my_array
	);
end entity;
-----------------------------------------------
architecture behavioral of CUTs is

	signal	w_Error	:	my_array(0 to g_N_Segments - 1)(g_N_Parallel - 1 downto 0) := (others => (others => '0'));

begin

	CUT_0:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(0));
	CUT_1:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(1));
	CUT_2:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(2));
	CUT_3:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(3));
	CUT_4:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(4));
	CUT_5:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(5));
	CUT_6:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(6));
	CUT_7:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(7));
	CUT_8:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(8));
	CUT_9:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(9));
	CUT_10:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(10));
	CUT_11:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(11));
	CUT_12:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(12));
	CUT_13:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(13));
	CUT_14:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(14));
	CUT_15:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(15));
	CUT_16:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(16));
	CUT_17:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(17));
	CUT_18:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(18));
	CUT_19:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(19));
	CUT_20:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(20));
	CUT_21:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(21));
	CUT_22:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(22));
	CUT_23:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(23));
	CUT_24:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(24));
	CUT_25:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(25));
	CUT_26:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(26));
	CUT_27:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(27));
	CUT_28:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(28));
	CUT_29:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(29));
	CUT_30:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(30));
	CUT_31:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(31));
	CUT_32:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(32));
	CUT_33:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(33));
	CUT_34:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(34));
	CUT_35:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(35));
	CUT_36:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(36));
	CUT_37:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(37));
	CUT_38:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(38));
	CUT_39:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(39));
	CUT_40:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(40));
	CUT_41:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(41));
	CUT_42:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(42));
	CUT_43:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(43));
	CUT_44:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(44));
	CUT_45:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(45));
	CUT_46:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(46));
	CUT_47:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(47));
	CUT_48:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(48));
	CUT_49:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(0)(49));
	CUT_50:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(0));
	CUT_51:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(1));
	CUT_52:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(2));
	CUT_53:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(3));
	CUT_54:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(4));
	CUT_55:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(5));
	CUT_56:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(6));
	CUT_57:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(7));
	CUT_58:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(8));
	CUT_59:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(9));
	CUT_60:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(10));
	CUT_61:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(11));
	CUT_62:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(12));
	CUT_63:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(13));
	CUT_64:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(14));
	CUT_65:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(15));
	CUT_66:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(16));
	CUT_67:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(17));
	CUT_68:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(18));
	CUT_69:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(19));
	CUT_70:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(20));
	CUT_71:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(21));
	CUT_72:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(22));
	CUT_73:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(23));
	CUT_74:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(24));
	CUT_75:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(25));
	CUT_76:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(26));
	CUT_77:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(27));
	CUT_78:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(28));
	CUT_79:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(29));
	CUT_80:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(30));
	CUT_81:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(31));
	CUT_82:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(32));
	CUT_83:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(33));
	CUT_84:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(34));
	CUT_85:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(35));
	CUT_86:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(36));
	CUT_87:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(37));
	CUT_88:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(38));
	CUT_89:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(39));
	CUT_90:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(40));
	CUT_91:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(41));
	CUT_92:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(42));
	CUT_93:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(43));
	CUT_94:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(44));
	CUT_95:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(45));
	CUT_96:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(46));
	CUT_97:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(47));
	CUT_98:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(48));
	CUT_99:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(1)(49));
	CUT_100:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(0));
	CUT_101:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(1));
	CUT_102:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(2));
	CUT_103:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(3));
	CUT_104:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(4));
	CUT_105:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(5));
	CUT_106:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(6));
	CUT_107:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(7));
	CUT_108:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(8));
	CUT_109:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(9));
	CUT_110:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(10));
	CUT_111:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(11));
	CUT_112:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(12));
	CUT_113:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(13));
	CUT_114:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(14));
	CUT_115:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(15));
	CUT_116:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(16));
	CUT_117:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(17));
	CUT_118:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(18));
	CUT_119:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(19));
	CUT_120:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(20));
	CUT_121:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(21));
	CUT_122:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(22));
	CUT_123:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(23));
	CUT_124:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(24));
	CUT_125:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(25));
	CUT_126:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(26));
	CUT_127:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(27));
	CUT_128:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(28));
	CUT_129:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(29));
	CUT_130:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(30));
	CUT_131:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(31));
	CUT_132:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(32));
	CUT_133:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(33));
	CUT_134:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(34));
	CUT_135:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(35));
	CUT_136:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(36));
	CUT_137:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(37));
	CUT_138:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(38));
	CUT_139:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(39));
	CUT_140:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(40));
	CUT_141:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(41));
	CUT_142:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(42));
	CUT_143:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(43));
	CUT_144:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(44));
	CUT_145:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(45));
	CUT_146:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(46));
	CUT_147:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(47));
	CUT_148:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(48));
	CUT_149:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(2)(49));
	CUT_150:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(0));
	CUT_151:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(1));
	CUT_152:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(2));
	CUT_153:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(3));
	CUT_154:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(4));
	CUT_155:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(5));
	CUT_156:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(6));
	CUT_157:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(7));
	CUT_158:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(8));
	CUT_159:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(9));
	CUT_160:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(10));
	CUT_161:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(11));
	CUT_162:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(12));
	CUT_163:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(13));
	CUT_164:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(14));
	CUT_165:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(15));
	CUT_166:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(16));
	CUT_167:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(17));
	CUT_168:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(18));
	CUT_169:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(19));
	CUT_170:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(20));
	CUT_171:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(21));
	CUT_172:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(22));
	CUT_173:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(23));
	CUT_174:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(24));
	CUT_175:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(25));
	CUT_176:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(26));
	CUT_177:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(27));
	CUT_178:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(28));
	CUT_179:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(29));
	CUT_180:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(30));
	CUT_181:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(31));
	CUT_182:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(32));
	CUT_183:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(33));
	CUT_184:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(34));
	CUT_185:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(35));
	CUT_186:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(36));
	CUT_187:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(37));
	CUT_188:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(38));
	CUT_189:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(39));
	CUT_190:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(40));
	CUT_191:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(41));
	CUT_192:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(42));
	CUT_193:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(43));
	CUT_194:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(44));
	CUT_195:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(45));
	CUT_196:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(46));
	CUT_197:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(47));
	CUT_198:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(48));
	CUT_199:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(3)(49));
	CUT_200:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(0));
	CUT_201:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(1));
	CUT_202:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(2));
	CUT_203:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(3));
	CUT_204:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(4));
	CUT_205:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(5));
	CUT_206:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(6));
	CUT_207:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(7));
	CUT_208:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(8));
	CUT_209:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(9));
	CUT_210:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(10));
	CUT_211:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(11));
	CUT_212:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(12));
	CUT_213:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(13));
	CUT_214:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(14));
	CUT_215:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(15));
	CUT_216:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(16));
	CUT_217:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(17));
	CUT_218:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(18));
	CUT_219:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(19));
	CUT_220:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(20));
	CUT_221:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(21));
	CUT_222:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(22));
	CUT_223:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(23));
	CUT_224:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(24));
	CUT_225:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(25));
	CUT_226:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(26));
	CUT_227:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(27));
	CUT_228:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(28));
	CUT_229:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(29));
	CUT_230:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(30));
	CUT_231:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(31));
	CUT_232:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(32));
	CUT_233:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(33));
	CUT_234:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(34));
	CUT_235:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(35));
	CUT_236:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(36));
	CUT_237:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(37));
	CUT_238:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(38));
	CUT_239:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(39));
	CUT_240:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(40));
	CUT_241:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(41));
	CUT_242:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(42));
	CUT_243:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(43));
	CUT_244:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(44));
	CUT_245:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(45));
	CUT_246:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(46));
	CUT_247:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(47));
	CUT_248:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(48));
	CUT_249:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(4)(49));
	CUT_250:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(0));
	CUT_251:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(1));
	CUT_252:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(2));
	CUT_253:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(3));
	CUT_254:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(4));
	CUT_255:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(5));
	CUT_256:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(6));
	CUT_257:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(7));
	CUT_258:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(8));
	CUT_259:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(9));
	CUT_260:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(10));
	CUT_261:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(11));
	CUT_262:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(12));
	CUT_263:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(13));
	CUT_264:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(14));
	CUT_265:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(15));
	CUT_266:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(16));
	CUT_267:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(17));
	CUT_268:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(18));
	CUT_269:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(19));
	CUT_270:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(20));
	CUT_271:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(21));
	CUT_272:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(22));
	CUT_273:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(23));
	CUT_274:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(24));
	CUT_275:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(25));
	CUT_276:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(26));
	CUT_277:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(27));
	CUT_278:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(28));
	CUT_279:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(29));
	CUT_280:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(30));
	CUT_281:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(31));
	CUT_282:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(32));
	CUT_283:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(33));
	CUT_284:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(34));
	CUT_285:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(35));
	CUT_286:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(36));
	CUT_287:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(37));
	CUT_288:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(38));
	CUT_289:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(39));
	CUT_290:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(40));
	CUT_291:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(41));
	CUT_292:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(42));
	CUT_293:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(43));
	CUT_294:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(44));
	CUT_295:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(45));
	CUT_296:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(46));
	CUT_297:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(47));
	CUT_298:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(48));
	CUT_299:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(5)(49));
	CUT_300:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(0));
	CUT_301:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(1));
	CUT_302:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(2));
	CUT_303:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(3));
	CUT_304:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(4));
	CUT_305:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(5));
	CUT_306:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(6));
	CUT_307:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(7));
	CUT_308:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(8));
	CUT_309:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(9));
	CUT_310:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(10));
	CUT_311:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(11));
	CUT_312:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(12));
	CUT_313:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(13));
	CUT_314:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(14));
	CUT_315:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(15));
	CUT_316:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(16));
	CUT_317:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(17));
	CUT_318:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(18));
	CUT_319:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(19));
	CUT_320:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(20));
	CUT_321:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(21));
	CUT_322:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(22));
	CUT_323:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(23));
	CUT_324:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(24));
	CUT_325:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(25));
	CUT_326:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(26));
	CUT_327:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(27));
	CUT_328:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(28));
	CUT_329:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(29));
	CUT_330:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(30));
	CUT_331:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(31));
	CUT_332:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(32));
	CUT_333:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(33));
	CUT_334:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(34));
	CUT_335:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(35));
	CUT_336:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(36));
	CUT_337:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(37));
	CUT_338:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(38));
	CUT_339:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(39));
	CUT_340:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(40));
	CUT_341:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(41));
	CUT_342:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(42));
	CUT_343:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(43));
	CUT_344:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(44));
	CUT_345:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(45));
	CUT_346:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(46));
	CUT_347:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(47));
	CUT_348:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(48));
	CUT_349:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(6)(49));
	CUT_350:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(0));
	CUT_351:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(1));
	CUT_352:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(2));
	CUT_353:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(3));
	CUT_354:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(4));
	CUT_355:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(5));
	CUT_356:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(6));
	CUT_357:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(7));
	CUT_358:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(8));
	CUT_359:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(9));
	CUT_360:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(10));
	CUT_361:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(11));
	CUT_362:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(12));
	CUT_363:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(13));
	CUT_364:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(14));
	CUT_365:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(15));
	CUT_366:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(16));
	CUT_367:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(17));
	CUT_368:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(18));
	CUT_369:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(19));
	CUT_370:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(20));
	CUT_371:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(21));
	CUT_372:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(22));
	CUT_373:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(23));
	CUT_374:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(24));
	CUT_375:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(25));
	CUT_376:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(26));
	CUT_377:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(27));
	CUT_378:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(28));
	CUT_379:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(29));
	CUT_380:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(30));
	CUT_381:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(31));
	CUT_382:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(32));
	CUT_383:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(33));
	CUT_384:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(34));
	CUT_385:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(35));
	CUT_386:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(36));
	CUT_387:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(37));
	CUT_388:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(38));
	CUT_389:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(39));
	CUT_390:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(40));
	CUT_391:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(41));
	CUT_392:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(42));
	CUT_393:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(43));
	CUT_394:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(44));
	CUT_395:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(45));
	CUT_396:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(46));
	CUT_397:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(47));
	CUT_398:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(48));
	CUT_399:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(7)(49));
	CUT_400:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(0));
	CUT_401:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(1));
	CUT_402:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(2));
	CUT_403:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(3));
	CUT_404:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(4));
	CUT_405:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(5));
	CUT_406:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(6));
	CUT_407:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(7));
	CUT_408:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(8));
	CUT_409:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(9));
	CUT_410:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(10));
	CUT_411:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(11));
	CUT_412:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(12));
	CUT_413:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(13));
	CUT_414:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(14));
	CUT_415:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(15));
	CUT_416:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(16));
	CUT_417:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(17));
	CUT_418:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(18));
	CUT_419:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(19));
	CUT_420:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(20));
	CUT_421:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(21));
	CUT_422:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(22));
	CUT_423:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(23));
	CUT_424:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(24));
	CUT_425:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(25));
	CUT_426:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(26));
	CUT_427:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(27));
	CUT_428:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(28));
	CUT_429:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(29));
	CUT_430:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(30));
	CUT_431:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(31));
	CUT_432:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(32));
	CUT_433:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(33));
	CUT_434:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(34));
	CUT_435:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(35));
	CUT_436:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(36));
	CUT_437:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(37));
	CUT_438:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(38));
	CUT_439:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(39));
	CUT_440:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(40));
	CUT_441:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(41));
	CUT_442:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(42));
	CUT_443:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(43));
	CUT_444:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(44));
	CUT_445:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(45));
	CUT_446:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(46));
	CUT_447:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(47));
	CUT_448:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(48));
	CUT_449:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(8)(49));
	CUT_450:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(0));
	CUT_451:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(1));
	CUT_452:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(2));
	CUT_453:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(3));
	CUT_454:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(4));
	CUT_455:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(5));
	CUT_456:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(6));
	CUT_457:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(7));
	CUT_458:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(8));
	CUT_459:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(9));
	CUT_460:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(10));
	CUT_461:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(11));
	CUT_462:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(12));
	CUT_463:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(13));
	CUT_464:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(14));
	CUT_465:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(15));
	CUT_466:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(16));
	CUT_467:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(17));
	CUT_468:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(18));
	CUT_469:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(19));
	CUT_470:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(20));
	CUT_471:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(21));
	CUT_472:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(22));
	CUT_473:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(23));
	CUT_474:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(24));
	CUT_475:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(25));
	CUT_476:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(26));
	CUT_477:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(27));
	CUT_478:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(28));
	CUT_479:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(29));
	CUT_480:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(30));
	CUT_481:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(31));
	CUT_482:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(32));
	CUT_483:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(33));
	CUT_484:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(34));
	CUT_485:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(35));
	CUT_486:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(36));
	CUT_487:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(37));
	CUT_488:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(38));
	CUT_489:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(39));
	CUT_490:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(40));
	CUT_491:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(41));
	CUT_492:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(42));
	CUT_493:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(43));
	CUT_494:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(44));
	CUT_495:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(45));
	CUT_496:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(46));
	CUT_497:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(47));
	CUT_498:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(48));
	CUT_499:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(9)(49));
	CUT_500:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(0));
	CUT_501:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(1));
	CUT_502:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(2));
	CUT_503:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(3));
	CUT_504:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(4));
	CUT_505:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(5));
	CUT_506:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(6));
	CUT_507:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(7));
	CUT_508:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(8));
	CUT_509:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(9));
	CUT_510:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(10));
	CUT_511:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(11));
	CUT_512:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(12));
	CUT_513:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(13));
	CUT_514:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(14));
	CUT_515:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(15));
	CUT_516:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(16));
	CUT_517:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(17));
	CUT_518:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(18));
	CUT_519:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(19));
	CUT_520:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(20));
	CUT_521:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(21));
	CUT_522:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(22));
	CUT_523:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(23));
	CUT_524:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(24));
	CUT_525:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(25));
	CUT_526:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(26));
	CUT_527:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(27));
	CUT_528:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(28));
	CUT_529:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(29));
	CUT_530:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(30));
	CUT_531:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(31));
	CUT_532:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(32));
	CUT_533:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(33));
	CUT_534:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(34));
	CUT_535:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(35));
	CUT_536:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(36));
	CUT_537:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(37));
	CUT_538:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(38));
	CUT_539:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(39));
	CUT_540:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(40));
	CUT_541:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(41));
	CUT_542:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(42));
	CUT_543:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(43));
	CUT_544:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(44));
	CUT_545:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(45));
	CUT_546:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(46));
	CUT_547:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(47));
	CUT_548:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(48));
	CUT_549:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(10)(49));
	CUT_550:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(0));
	CUT_551:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(1));
	CUT_552:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(2));
	CUT_553:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(3));
	CUT_554:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(4));
	CUT_555:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(5));
	CUT_556:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(6));
	CUT_557:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(7));
	CUT_558:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(8));
	CUT_559:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(9));
	CUT_560:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(10));
	CUT_561:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(11));
	CUT_562:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(12));
	CUT_563:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(13));
	CUT_564:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(14));
	CUT_565:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(15));
	CUT_566:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(16));
	CUT_567:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(17));
	CUT_568:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(18));
	CUT_569:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(19));
	CUT_570:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(20));
	CUT_571:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(21));
	CUT_572:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(22));
	CUT_573:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(23));
	CUT_574:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(24));
	CUT_575:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(25));
	CUT_576:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(26));
	CUT_577:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(27));
	CUT_578:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(28));
	CUT_579:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(29));
	CUT_580:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(30));
	CUT_581:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(31));
	CUT_582:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(32));
	CUT_583:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(33));
	CUT_584:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(34));
	CUT_585:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(35));
	CUT_586:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(36));
	CUT_587:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(37));
	CUT_588:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(38));
	CUT_589:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(39));
	CUT_590:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(40));
	CUT_591:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(41));
	CUT_592:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(42));
	CUT_593:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(43));
	CUT_594:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(44));
	CUT_595:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(45));
	CUT_596:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(46));
	CUT_597:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(47));
	CUT_598:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(48));
	CUT_599:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(11)(49));
	CUT_600:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(0));
	CUT_601:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(1));
	CUT_602:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(2));
	CUT_603:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(3));
	CUT_604:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(4));
	CUT_605:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(5));
	CUT_606:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(6));
	CUT_607:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(7));
	CUT_608:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(8));
	CUT_609:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(9));
	CUT_610:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(10));
	CUT_611:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(11));
	CUT_612:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(12));
	CUT_613:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(13));
	CUT_614:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(14));
	CUT_615:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(15));
	CUT_616:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(16));
	CUT_617:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(17));
	CUT_618:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(18));
	CUT_619:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(19));
	CUT_620:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(20));
	CUT_621:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(21));
	CUT_622:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(22));
	CUT_623:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(23));
	CUT_624:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(24));
	CUT_625:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(25));
	CUT_626:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(26));
	CUT_627:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(27));
	CUT_628:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(28));
	CUT_629:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(29));
	CUT_630:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(30));
	CUT_631:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(31));
	CUT_632:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(32));
	CUT_633:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(33));
	CUT_634:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(34));
	CUT_635:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(35));
	CUT_636:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(36));
	CUT_637:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(37));
	CUT_638:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(38));
	CUT_639:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(39));
	CUT_640:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(40));
	CUT_641:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(41));
	CUT_642:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(42));
	CUT_643:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(43));
	CUT_644:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(44));
	CUT_645:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(45));
	CUT_646:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(46));
	CUT_647:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(47));
	CUT_648:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(48));
	CUT_649:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(12)(49));
	CUT_650:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(0));
	CUT_651:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(1));
	CUT_652:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(2));
	CUT_653:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(3));
	CUT_654:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(4));
	CUT_655:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(5));
	CUT_656:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(6));
	CUT_657:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(7));
	CUT_658:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(8));
	CUT_659:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(9));
	CUT_660:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(10));
	CUT_661:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(11));
	CUT_662:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(12));
	CUT_663:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(13));
	CUT_664:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(14));
	CUT_665:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(15));
	CUT_666:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(16));
	CUT_667:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(17));
	CUT_668:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(18));
	CUT_669:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(19));
	CUT_670:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(20));
	CUT_671:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(21));
	CUT_672:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(22));
	CUT_673:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(23));
	CUT_674:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(24));
	CUT_675:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(25));
	CUT_676:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(26));
	CUT_677:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(27));
	CUT_678:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(28));
	CUT_679:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(29));
	CUT_680:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(30));
	CUT_681:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(31));
	CUT_682:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(32));
	CUT_683:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(33));
	CUT_684:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(34));
	CUT_685:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(35));
	CUT_686:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(36));
	CUT_687:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(37));
	CUT_688:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(38));
	CUT_689:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(39));
	CUT_690:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(40));
	CUT_691:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(41));
	CUT_692:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(42));
	CUT_693:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(43));
	CUT_694:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(44));
	CUT_695:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(45));
	CUT_696:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(46));
	CUT_697:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(47));
	CUT_698:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(48));
	CUT_699:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(13)(49));
	CUT_700:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(0));
	CUT_701:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(1));
	CUT_702:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(2));
	CUT_703:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(3));
	CUT_704:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(4));
	CUT_705:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(5));
	CUT_706:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(6));
	CUT_707:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(7));
	CUT_708:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(8));
	CUT_709:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(9));
	CUT_710:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(10));
	CUT_711:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(11));
	CUT_712:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(12));
	CUT_713:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(13));
	CUT_714:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(14));
	CUT_715:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(15));
	CUT_716:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(16));
	CUT_717:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(17));
	CUT_718:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(18));
	CUT_719:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(19));
	CUT_720:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(20));
	CUT_721:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(21));
	CUT_722:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(22));
	CUT_723:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(23));
	CUT_724:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(24));
	CUT_725:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(25));
	CUT_726:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(26));
	CUT_727:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(27));
	CUT_728:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(28));
	CUT_729:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(29));
	CUT_730:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(30));
	CUT_731:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(31));
	CUT_732:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(32));
	CUT_733:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(33));
	CUT_734:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(34));
	CUT_735:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(35));
	CUT_736:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(36));
	CUT_737:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(37));
	CUT_738:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(38));
	CUT_739:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(39));
	CUT_740:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(40));
	CUT_741:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(41));
	CUT_742:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(42));
	CUT_743:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(43));
	CUT_744:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(44));
	CUT_745:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(45));
	CUT_746:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(46));
	CUT_747:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(47));
	CUT_748:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(48));
	CUT_749:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(14)(49));
	CUT_750:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(0));
	CUT_751:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(1));
	CUT_752:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(2));
	CUT_753:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(3));
	CUT_754:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(4));
	CUT_755:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(5));
	CUT_756:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(6));
	CUT_757:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(7));
	CUT_758:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(8));
	CUT_759:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(9));
	CUT_760:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(10));
	CUT_761:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(11));
	CUT_762:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(12));
	CUT_763:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(13));
	CUT_764:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(14));
	CUT_765:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(15));
	CUT_766:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(16));
	CUT_767:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(17));
	CUT_768:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(18));
	CUT_769:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(19));
	CUT_770:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(20));
	CUT_771:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(21));
	CUT_772:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(22));
	CUT_773:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(23));
	CUT_774:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(24));
	CUT_775:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(25));
	CUT_776:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(26));
	CUT_777:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(27));
	CUT_778:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(28));
	CUT_779:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(29));
	CUT_780:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(30));
	CUT_781:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(31));
	CUT_782:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(32));
	CUT_783:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(33));
	CUT_784:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(34));
	CUT_785:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(35));
	CUT_786:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(36));
	CUT_787:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(37));
	CUT_788:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(38));
	CUT_789:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(39));
	CUT_790:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(40));
	CUT_791:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(41));
	CUT_792:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(42));
	CUT_793:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(43));
	CUT_794:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(44));
	CUT_795:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(45));
	CUT_796:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(46));
	CUT_797:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(47));
	CUT_798:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(48));
	CUT_799:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(15)(49));
	CUT_800:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(0));
	CUT_801:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(1));
	CUT_802:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(2));
	CUT_803:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(3));
	CUT_804:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(4));
	CUT_805:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(5));
	CUT_806:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(6));
	CUT_807:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(7));
	CUT_808:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(8));
	CUT_809:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(9));
	CUT_810:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(10));
	CUT_811:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(11));
	CUT_812:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(12));
	CUT_813:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(13));
	CUT_814:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(14));
	CUT_815:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(15));
	CUT_816:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(16));
	CUT_817:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(17));
	CUT_818:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(18));
	CUT_819:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(19));
	CUT_820:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(20));
	CUT_821:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(21));
	CUT_822:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(22));
	CUT_823:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(23));
	CUT_824:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(24));
	CUT_825:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(25));
	CUT_826:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(26));
	CUT_827:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(27));
	CUT_828:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(28));
	CUT_829:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(29));
	CUT_830:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(30));
	CUT_831:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(31));
	CUT_832:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(32));
	CUT_833:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(33));
	CUT_834:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(34));
	CUT_835:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(35));
	CUT_836:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(36));
	CUT_837:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(37));
	CUT_838:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(38));
	CUT_839:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(39));
	CUT_840:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(40));
	CUT_841:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(41));
	CUT_842:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(42));
	CUT_843:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(43));
	CUT_844:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(44));
	CUT_845:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(45));
	CUT_846:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(46));
	CUT_847:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(47));
	CUT_848:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(48));
	CUT_849:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(16)(49));
	CUT_850:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(0));
	CUT_851:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(1));
	CUT_852:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(2));
	CUT_853:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(3));
	CUT_854:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(4));
	CUT_855:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(5));
	CUT_856:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(6));
	CUT_857:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(7));
	CUT_858:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(8));
	CUT_859:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(9));
	CUT_860:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(10));
	CUT_861:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(11));
	CUT_862:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(12));
	CUT_863:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(13));
	CUT_864:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(14));
	CUT_865:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(15));
	CUT_866:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(16));
	CUT_867:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(17));
	CUT_868:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(18));
	CUT_869:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(19));
	CUT_870:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(20));
	CUT_871:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(21));
	CUT_872:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(22));
	CUT_873:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(23));
	CUT_874:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(24));
	CUT_875:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(25));
	CUT_876:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(26));
	CUT_877:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(27));
	CUT_878:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(28));
	CUT_879:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(29));
	CUT_880:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(30));
	CUT_881:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(31));
	CUT_882:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(32));
	CUT_883:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(33));
	CUT_884:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(34));
	CUT_885:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(35));
	CUT_886:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(36));
	CUT_887:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(37));
	CUT_888:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(38));
	CUT_889:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(39));
	CUT_890:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(40));
	CUT_891:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(41));
	CUT_892:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(42));
	CUT_893:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(43));
	CUT_894:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(44));
	CUT_895:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(45));
	CUT_896:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(46));
	CUT_897:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(47));
	CUT_898:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(48));
	CUT_899:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(17)(49));
	CUT_900:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(0));
	CUT_901:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(1));
	CUT_902:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(2));
	CUT_903:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(3));
	CUT_904:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(4));
	CUT_905:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(5));
	CUT_906:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(6));
	CUT_907:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(7));
	CUT_908:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(8));
	CUT_909:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(9));
	CUT_910:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(10));
	CUT_911:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(11));
	CUT_912:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(12));
	CUT_913:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(13));
	CUT_914:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(14));
	CUT_915:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(15));
	CUT_916:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(16));
	CUT_917:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(17));
	CUT_918:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(18));
	CUT_919:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(19));
	CUT_920:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(20));
	CUT_921:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(21));
	CUT_922:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(22));
	CUT_923:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(23));
	CUT_924:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(24));
	CUT_925:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(25));
	CUT_926:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(26));
	CUT_927:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(27));
	CUT_928:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(28));
	CUT_929:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(29));
	CUT_930:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(30));
	CUT_931:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(31));
	CUT_932:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(32));
	CUT_933:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(33));
	CUT_934:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(34));
	CUT_935:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(35));
	CUT_936:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(36));
	CUT_937:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(37));
	CUT_938:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(38));
	CUT_939:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(39));
	CUT_940:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(40));
	CUT_941:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(41));
	CUT_942:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(42));
	CUT_943:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(43));
	CUT_944:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(44));
	CUT_945:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(45));
	CUT_946:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(46));
	CUT_947:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(47));
	CUT_948:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(48));
	CUT_949:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(18)(49));
	CUT_950:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(0));
	CUT_951:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(1));
	CUT_952:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(2));
	CUT_953:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(3));
	CUT_954:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(4));
	CUT_955:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(5));
	CUT_956:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(6));
	CUT_957:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(7));
	CUT_958:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(8));
	CUT_959:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(9));
	CUT_960:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(10));
	CUT_961:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(11));
	CUT_962:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(12));
	CUT_963:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(13));
	CUT_964:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(14));
	CUT_965:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(15));
	CUT_966:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(16));
	CUT_967:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(17));
	CUT_968:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(18));
	CUT_969:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(19));
	CUT_970:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(20));
	CUT_971:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(21));
	CUT_972:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(22));
	CUT_973:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(23));
	CUT_974:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(24));
	CUT_975:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(25));
	CUT_976:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(26));
	CUT_977:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(27));
	CUT_978:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(28));
	CUT_979:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(29));
	CUT_980:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(30));
	CUT_981:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(31));
	CUT_982:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(32));
	CUT_983:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(33));
	CUT_984:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(34));
	CUT_985:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(35));
	CUT_986:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(36));
	CUT_987:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(37));
	CUT_988:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(38));
	CUT_989:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(39));
	CUT_990:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(40));
	CUT_991:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(41));
	CUT_992:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(42));
	CUT_993:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(43));
	CUT_994:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(44));
	CUT_995:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(45));
	CUT_996:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(46));
	CUT_997:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(47));
	CUT_998:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(48));
	CUT_999:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(19)(49));
	CUT_1000:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(0));
	CUT_1001:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(1));
	CUT_1002:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(2));
	CUT_1003:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(3));
	CUT_1004:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(4));
	CUT_1005:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(5));
	CUT_1006:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(6));
	CUT_1007:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(7));
	CUT_1008:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(8));
	CUT_1009:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(9));
	CUT_1010:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(10));
	CUT_1011:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(11));
	CUT_1012:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(12));
	CUT_1013:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(13));
	CUT_1014:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(14));
	CUT_1015:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(15));
	CUT_1016:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(16));
	CUT_1017:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(17));
	CUT_1018:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(18));
	CUT_1019:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(19));
	CUT_1020:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(20));
	CUT_1021:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(21));
	CUT_1022:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(22));
	CUT_1023:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(23));
	CUT_1024:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(24));
	CUT_1025:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(25));
	CUT_1026:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(26));
	CUT_1027:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(27));
	CUT_1028:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(28));
	CUT_1029:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(29));
	CUT_1030:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(30));
	CUT_1031:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(31));
	CUT_1032:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(32));
	CUT_1033:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(33));
	CUT_1034:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(34));
	CUT_1035:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(35));
	CUT_1036:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(36));
	CUT_1037:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(37));
	CUT_1038:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(38));
	CUT_1039:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(39));
	CUT_1040:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(40));
	CUT_1041:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(41));
	CUT_1042:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(42));
	CUT_1043:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(43));
	CUT_1044:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(44));
	CUT_1045:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(45));
	CUT_1046:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(46));
	CUT_1047:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(47));
	CUT_1048:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(48));
	CUT_1049:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(20)(49));
	CUT_1050:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(0));
	CUT_1051:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(1));
	CUT_1052:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(2));
	CUT_1053:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(3));
	CUT_1054:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(4));
	CUT_1055:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(5));
	CUT_1056:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(6));
	CUT_1057:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(7));
	CUT_1058:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(8));
	CUT_1059:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(9));
	CUT_1060:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(10));
	CUT_1061:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(11));
	CUT_1062:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(12));
	CUT_1063:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(13));
	CUT_1064:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(14));
	CUT_1065:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(15));
	CUT_1066:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(16));
	CUT_1067:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(17));
	CUT_1068:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(18));
	CUT_1069:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(19));
	CUT_1070:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(20));
	CUT_1071:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(21));
	CUT_1072:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(22));
	CUT_1073:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(23));
	CUT_1074:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(24));
	CUT_1075:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(25));
	CUT_1076:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(26));
	CUT_1077:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(27));
	CUT_1078:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(28));
	CUT_1079:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(29));
	CUT_1080:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(30));
	CUT_1081:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(31));
	CUT_1082:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(32));
	CUT_1083:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(33));
	CUT_1084:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(34));
	CUT_1085:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(35));
	CUT_1086:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(36));
	CUT_1087:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(37));
	CUT_1088:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(38));
	CUT_1089:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(39));
	CUT_1090:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(40));
	CUT_1091:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(41));
	CUT_1092:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(42));
	CUT_1093:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(43));
	CUT_1094:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(44));
	CUT_1095:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(45));
	CUT_1096:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(46));
	CUT_1097:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(47));
	CUT_1098:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(48));
	CUT_1099:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(21)(49));
	CUT_1100:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(0));
	CUT_1101:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(1));
	CUT_1102:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(2));
	CUT_1103:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(3));
	CUT_1104:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(4));
	CUT_1105:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(5));
	CUT_1106:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(6));
	CUT_1107:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(7));
	CUT_1108:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(8));
	CUT_1109:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(9));
	CUT_1110:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(10));
	CUT_1111:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(11));
	CUT_1112:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(12));
	CUT_1113:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(13));
	CUT_1114:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(14));
	CUT_1115:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(15));
	CUT_1116:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(16));
	CUT_1117:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(17));
	CUT_1118:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(18));
	CUT_1119:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(19));
	CUT_1120:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(20));
	CUT_1121:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(21));
	CUT_1122:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(22));
	CUT_1123:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(23));
	CUT_1124:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(24));
	CUT_1125:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(25));
	CUT_1126:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(26));
	CUT_1127:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(27));
	CUT_1128:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(28));
	CUT_1129:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(29));
	CUT_1130:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(30));
	CUT_1131:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(31));
	CUT_1132:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(32));
	CUT_1133:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(33));
	CUT_1134:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(34));
	CUT_1135:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(35));
	CUT_1136:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(36));
	CUT_1137:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(37));
	CUT_1138:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(38));
	CUT_1139:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(39));
	CUT_1140:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(40));
	CUT_1141:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(41));
	CUT_1142:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(42));
	CUT_1143:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(43));
	CUT_1144:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(44));
	CUT_1145:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(45));
	CUT_1146:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(46));
	CUT_1147:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(47));
	CUT_1148:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(48));
	CUT_1149:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(22)(49));
	CUT_1150:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(0));
	CUT_1151:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(1));
	CUT_1152:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(2));
	CUT_1153:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(3));
	CUT_1154:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(4));
	CUT_1155:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(5));
	CUT_1156:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(6));
	CUT_1157:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(7));
	CUT_1158:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(8));
	CUT_1159:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(9));
	CUT_1160:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(10));
	CUT_1161:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(11));
	CUT_1162:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(12));
	CUT_1163:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(13));
	CUT_1164:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(14));
	CUT_1165:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(15));
	CUT_1166:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(16));
	CUT_1167:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(17));
	CUT_1168:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(18));
	CUT_1169:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(19));
	CUT_1170:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(20));
	CUT_1171:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(21));
	CUT_1172:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(22));
	CUT_1173:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(23));
	CUT_1174:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(24));
	CUT_1175:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(25));
	CUT_1176:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(26));
	CUT_1177:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(27));
	CUT_1178:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(28));
	CUT_1179:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(29));
	CUT_1180:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(30));
	CUT_1181:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(31));
	CUT_1182:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(32));
	CUT_1183:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(33));
	CUT_1184:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(34));
	CUT_1185:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(35));
	CUT_1186:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(36));
	CUT_1187:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(37));
	CUT_1188:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(38));
	CUT_1189:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(39));
	CUT_1190:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(40));
	CUT_1191:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(41));
	CUT_1192:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(42));
	CUT_1193:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(43));
	CUT_1194:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(44));
	CUT_1195:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(45));
	CUT_1196:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(46));
	CUT_1197:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(47));
	CUT_1198:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(48));
	CUT_1199:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(23)(49));
	CUT_1200:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(0));
	CUT_1201:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(1));
	CUT_1202:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(2));
	CUT_1203:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(3));
	CUT_1204:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(4));
	CUT_1205:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(5));
	CUT_1206:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(6));
	CUT_1207:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(7));
	CUT_1208:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(8));
	CUT_1209:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(9));
	CUT_1210:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(10));
	CUT_1211:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(11));
	CUT_1212:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(12));
	CUT_1213:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(13));
	CUT_1214:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(14));
	CUT_1215:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(15));
	CUT_1216:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(16));
	CUT_1217:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(17));
	CUT_1218:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(18));
	CUT_1219:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(19));
	CUT_1220:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(20));
	CUT_1221:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(21));
	CUT_1222:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(22));
	CUT_1223:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(23));
	CUT_1224:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(24));
	CUT_1225:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(25));
	CUT_1226:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(26));
	CUT_1227:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(27));
	CUT_1228:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(28));
	CUT_1229:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(29));
	CUT_1230:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(30));
	CUT_1231:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(31));
	CUT_1232:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(32));
	CUT_1233:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(33));
	CUT_1234:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(34));
	CUT_1235:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(35));
	CUT_1236:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(36));
	CUT_1237:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(37));
	CUT_1238:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(38));
	CUT_1239:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(39));
	CUT_1240:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(40));
	CUT_1241:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(41));
	CUT_1242:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(42));
	CUT_1243:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(43));
	CUT_1244:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(44));
	CUT_1245:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(45));
	CUT_1246:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(46));
	CUT_1247:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(47));
	CUT_1248:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(48));
	CUT_1249:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(24)(49));
	CUT_1250:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(0));
	CUT_1251:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(1));
	CUT_1252:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(2));
	CUT_1253:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(3));
	CUT_1254:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(4));
	CUT_1255:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(5));
	CUT_1256:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(6));
	CUT_1257:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(7));
	CUT_1258:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(8));
	CUT_1259:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(9));
	CUT_1260:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(10));
	CUT_1261:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(11));
	CUT_1262:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(12));
	CUT_1263:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(13));
	CUT_1264:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(14));
	CUT_1265:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(15));
	CUT_1266:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(16));
	CUT_1267:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(17));
	CUT_1268:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(18));
	CUT_1269:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(19));
	CUT_1270:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(20));
	CUT_1271:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(21));
	CUT_1272:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(22));
	CUT_1273:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(23));
	CUT_1274:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(24));
	CUT_1275:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(25));
	CUT_1276:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(26));
	CUT_1277:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(27));
	CUT_1278:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(28));
	CUT_1279:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(29));
	CUT_1280:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(30));
	CUT_1281:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(31));
	CUT_1282:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(32));
	CUT_1283:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(33));
	CUT_1284:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(34));
	CUT_1285:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(35));
	CUT_1286:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(36));
	CUT_1287:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(37));
	CUT_1288:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(38));
	CUT_1289:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(39));
	CUT_1290:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(40));
	CUT_1291:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(41));
	CUT_1292:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(42));
	CUT_1293:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(43));
	CUT_1294:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(44));
	CUT_1295:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(45));
	CUT_1296:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(46));
	CUT_1297:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(47));
	CUT_1298:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(48));
	CUT_1299:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(25)(49));
	CUT_1300:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(0));
	CUT_1301:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(1));
	CUT_1302:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(2));
	CUT_1303:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(3));
	CUT_1304:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(4));
	CUT_1305:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(5));
	CUT_1306:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(6));
	CUT_1307:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(7));
	CUT_1308:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(8));
	CUT_1309:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(9));
	CUT_1310:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(10));
	CUT_1311:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(11));
	CUT_1312:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(12));
	CUT_1313:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(13));
	CUT_1314:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(14));
	CUT_1315:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(15));
	CUT_1316:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(16));
	CUT_1317:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(17));
	CUT_1318:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(18));
	CUT_1319:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(19));
	CUT_1320:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(20));
	CUT_1321:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(21));
	CUT_1322:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(22));
	CUT_1323:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(23));
	CUT_1324:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(24));
	CUT_1325:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(25));
	CUT_1326:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(26));
	CUT_1327:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(27));
	CUT_1328:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(28));
	CUT_1329:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(29));
	CUT_1330:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(30));
	CUT_1331:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(31));
	CUT_1332:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(32));
	CUT_1333:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(33));
	CUT_1334:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(34));
	CUT_1335:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(35));
	CUT_1336:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(36));
	CUT_1337:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(37));
	CUT_1338:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(38));
	CUT_1339:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(39));
	CUT_1340:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(40));
	CUT_1341:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(41));
	CUT_1342:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(42));
	CUT_1343:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(43));
	CUT_1344:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(44));
	CUT_1345:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(45));
	CUT_1346:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(46));
	CUT_1347:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(47));
	CUT_1348:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(48));
	CUT_1349:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(26)(49));
	CUT_1350:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(0));
	CUT_1351:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(1));
	CUT_1352:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(2));
	CUT_1353:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(3));
	CUT_1354:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(4));
	CUT_1355:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(5));
	CUT_1356:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(6));
	CUT_1357:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(7));
	CUT_1358:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(8));
	CUT_1359:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(9));
	CUT_1360:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(10));
	CUT_1361:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(11));
	CUT_1362:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(12));
	CUT_1363:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(13));
	CUT_1364:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(14));
	CUT_1365:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(15));
	CUT_1366:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(16));
	CUT_1367:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(17));
	CUT_1368:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(18));
	CUT_1369:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(19));
	CUT_1370:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(20));
	CUT_1371:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(21));
	CUT_1372:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(22));
	CUT_1373:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(23));
	CUT_1374:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(24));
	CUT_1375:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(25));
	CUT_1376:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(26));
	CUT_1377:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(27));
	CUT_1378:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(28));
	CUT_1379:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(29));
	CUT_1380:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(30));
	CUT_1381:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(31));
	CUT_1382:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(32));
	CUT_1383:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(33));
	CUT_1384:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(34));
	CUT_1385:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(35));
	CUT_1386:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(36));
	CUT_1387:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(37));
	CUT_1388:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(38));
	CUT_1389:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(39));
	CUT_1390:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(40));
	CUT_1391:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(41));
	CUT_1392:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(42));
	CUT_1393:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(43));
	CUT_1394:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(44));
	CUT_1395:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(45));
	CUT_1396:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(46));
	CUT_1397:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(47));
	CUT_1398:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(48));
	CUT_1399:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(27)(49));
	CUT_1400:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(0));
	CUT_1401:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(1));
	CUT_1402:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(2));
	CUT_1403:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(3));
	CUT_1404:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(4));
	CUT_1405:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(5));
	CUT_1406:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(6));
	CUT_1407:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(7));
	CUT_1408:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(8));
	CUT_1409:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(9));
	CUT_1410:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(10));
	CUT_1411:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(11));
	CUT_1412:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(12));
	CUT_1413:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(13));
	CUT_1414:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(14));
	CUT_1415:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(15));
	CUT_1416:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(16));
	CUT_1417:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(17));
	CUT_1418:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(18));
	CUT_1419:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(19));
	CUT_1420:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(20));
	CUT_1421:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(21));
	CUT_1422:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(22));
	CUT_1423:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(23));
	CUT_1424:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(24));
	CUT_1425:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(25));
	CUT_1426:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(26));
	CUT_1427:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(27));
	CUT_1428:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(28));
	CUT_1429:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(29));
	CUT_1430:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(30));
	CUT_1431:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(31));
	CUT_1432:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(32));
	CUT_1433:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(33));
	CUT_1434:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(34));
	CUT_1435:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(35));
	CUT_1436:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(36));
	CUT_1437:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(37));
	CUT_1438:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(38));
	CUT_1439:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(39));
	CUT_1440:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(40));
	CUT_1441:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(41));
	CUT_1442:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(42));
	CUT_1443:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(43));
	CUT_1444:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(44));
	CUT_1445:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(45));
	CUT_1446:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(46));
	CUT_1447:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(47));
	CUT_1448:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(48));
	CUT_1449:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(28)(49));
	CUT_1450:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(0));
	CUT_1451:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(1));
	CUT_1452:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(2));
	CUT_1453:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(3));
	CUT_1454:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(4));
	CUT_1455:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(5));
	CUT_1456:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(6));
	CUT_1457:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(7));
	CUT_1458:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(8));
	CUT_1459:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(9));
	CUT_1460:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(10));
	CUT_1461:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(11));
	CUT_1462:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(12));
	CUT_1463:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(13));
	CUT_1464:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(14));
	CUT_1465:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(15));
	CUT_1466:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(16));
	CUT_1467:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(17));
	CUT_1468:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(18));
	CUT_1469:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(19));
	CUT_1470:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(20));
	CUT_1471:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(21));
	CUT_1472:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(22));
	CUT_1473:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(23));
	CUT_1474:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(24));
	CUT_1475:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(25));
	CUT_1476:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(26));
	CUT_1477:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(27));
	CUT_1478:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(28));
	CUT_1479:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(29));
	CUT_1480:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(30));
	CUT_1481:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(31));
	CUT_1482:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(32));
	CUT_1483:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(33));
	CUT_1484:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(34));
	CUT_1485:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(35));
	CUT_1486:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(36));
	CUT_1487:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(37));
	CUT_1488:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(38));
	CUT_1489:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(39));
	CUT_1490:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(40));
	CUT_1491:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(41));
	CUT_1492:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(42));
	CUT_1493:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(43));
	CUT_1494:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(44));
	CUT_1495:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(45));
	CUT_1496:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(46));
	CUT_1497:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(47));
	CUT_1498:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(48));
	CUT_1499:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(29)(49));
	CUT_1500:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(0));
	CUT_1501:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(1));
	CUT_1502:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(2));
	CUT_1503:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(3));
	CUT_1504:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(4));
	CUT_1505:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(5));
	CUT_1506:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(6));
	CUT_1507:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(7));
	CUT_1508:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(8));
	CUT_1509:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(9));
	CUT_1510:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(10));
	CUT_1511:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(11));
	CUT_1512:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(12));
	CUT_1513:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(13));
	CUT_1514:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(14));
	CUT_1515:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(15));
	CUT_1516:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(16));
	CUT_1517:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(17));
	CUT_1518:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(18));
	CUT_1519:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(19));
	CUT_1520:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(20));
	CUT_1521:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(21));
	CUT_1522:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(22));
	CUT_1523:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(23));
	CUT_1524:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(24));
	CUT_1525:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(25));
	CUT_1526:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(26));
	CUT_1527:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(27));
	CUT_1528:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(28));
	CUT_1529:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(29));
	CUT_1530:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(30));
	CUT_1531:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(31));
	CUT_1532:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(32));
	CUT_1533:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(33));
	CUT_1534:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(34));
	CUT_1535:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(35));
	CUT_1536:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(36));
	CUT_1537:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(37));
	CUT_1538:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(38));
	CUT_1539:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(39));
	CUT_1540:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(40));
	CUT_1541:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(41));
	CUT_1542:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(42));
	CUT_1543:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(43));
	CUT_1544:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(44));
	CUT_1545:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(45));
	CUT_1546:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(46));
	CUT_1547:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(47));
	CUT_1548:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(48));
	CUT_1549:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(30)(49));
	CUT_1550:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(0));
	CUT_1551:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(1));
	CUT_1552:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(2));
	CUT_1553:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(3));
	CUT_1554:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(4));
	CUT_1555:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(5));
	CUT_1556:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(6));
	CUT_1557:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(7));
	CUT_1558:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(8));
	CUT_1559:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(9));
	CUT_1560:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(10));
	CUT_1561:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(11));
	CUT_1562:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(12));
	CUT_1563:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(13));
	CUT_1564:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(14));
	CUT_1565:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(15));
	CUT_1566:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(16));
	CUT_1567:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(17));
	CUT_1568:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(18));
	CUT_1569:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(19));
	CUT_1570:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(20));
	CUT_1571:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(21));
	CUT_1572:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(22));
	CUT_1573:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(23));
	CUT_1574:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(24));
	CUT_1575:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(25));
	CUT_1576:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(26));
	CUT_1577:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(27));
	CUT_1578:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(28));
	CUT_1579:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(29));
	CUT_1580:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(30));
	CUT_1581:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(31));
	CUT_1582:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(32));
	CUT_1583:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(33));
	CUT_1584:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(34));
	CUT_1585:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(35));
	CUT_1586:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(36));
	CUT_1587:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(37));
	CUT_1588:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(38));
	CUT_1589:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(39));
	CUT_1590:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(40));
	CUT_1591:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(41));
	CUT_1592:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(42));
	CUT_1593:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(43));
	CUT_1594:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(44));
	CUT_1595:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(45));
	CUT_1596:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(46));
	CUT_1597:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(47));
	CUT_1598:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(48));
	CUT_1599:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(31)(49));
	CUT_1600:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(0));
	CUT_1601:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(1));
	CUT_1602:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(2));
	CUT_1603:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(3));
	CUT_1604:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(4));
	CUT_1605:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(5));
	CUT_1606:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(6));
	CUT_1607:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(7));
	CUT_1608:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(8));
	CUT_1609:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(9));
	CUT_1610:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(10));
	CUT_1611:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(11));
	CUT_1612:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(12));
	CUT_1613:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(13));
	CUT_1614:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(14));
	CUT_1615:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(15));
	CUT_1616:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(16));
	CUT_1617:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(17));
	CUT_1618:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(18));
	CUT_1619:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(19));
	CUT_1620:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(20));
	CUT_1621:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(21));
	CUT_1622:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(22));
	CUT_1623:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(23));
	CUT_1624:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(24));
	CUT_1625:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(25));
	CUT_1626:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(26));
	CUT_1627:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(27));
	CUT_1628:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(28));
	CUT_1629:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(29));
	CUT_1630:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(30));
	CUT_1631:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(31));
	CUT_1632:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(32));
	CUT_1633:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(33));
	CUT_1634:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(34));
	CUT_1635:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(35));
	CUT_1636:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(36));
	CUT_1637:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(37));
	CUT_1638:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(38));
	CUT_1639:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(39));
	CUT_1640:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(40));
	CUT_1641:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(41));
	CUT_1642:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(42));
	CUT_1643:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(43));
	CUT_1644:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(44));
	CUT_1645:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(45));
	CUT_1646:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(46));
	CUT_1647:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(47));
	CUT_1648:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(48));
	CUT_1649:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(32)(49));
	CUT_1650:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(0));
	CUT_1651:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(1));
	CUT_1652:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(2));
	CUT_1653:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(3));
	CUT_1654:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(4));
	CUT_1655:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(5));
	CUT_1656:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(6));
	CUT_1657:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(7));
	CUT_1658:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(8));
	CUT_1659:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(9));
	CUT_1660:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(10));
	CUT_1661:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(11));
	CUT_1662:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(12));
	CUT_1663:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(13));
	CUT_1664:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(14));
	CUT_1665:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(15));
	CUT_1666:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(16));
	CUT_1667:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(17));
	CUT_1668:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(18));
	CUT_1669:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(19));
	CUT_1670:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(20));
	CUT_1671:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(21));
	CUT_1672:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(22));
	CUT_1673:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(23));
	CUT_1674:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(24));
	CUT_1675:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(25));
	CUT_1676:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(26));
	CUT_1677:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(27));
	CUT_1678:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(28));
	CUT_1679:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(29));
	CUT_1680:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(30));
	CUT_1681:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(31));
	CUT_1682:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(32));
	CUT_1683:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(33));
	CUT_1684:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(34));
	CUT_1685:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(35));
	CUT_1686:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(36));
	CUT_1687:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(37));
	CUT_1688:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(38));
	CUT_1689:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(39));
	CUT_1690:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(40));
	CUT_1691:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(41));
	CUT_1692:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(42));
	CUT_1693:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(43));
	CUT_1694:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(44));
	CUT_1695:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(45));
	CUT_1696:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(46));
	CUT_1697:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(47));
	CUT_1698:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(48));
	CUT_1699:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(33)(49));
	CUT_1700:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(0));
	CUT_1701:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(1));
	CUT_1702:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(2));
	CUT_1703:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(3));
	CUT_1704:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(4));
	CUT_1705:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(5));
	CUT_1706:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(6));
	CUT_1707:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(7));
	CUT_1708:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(8));
	CUT_1709:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(9));
	CUT_1710:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(10));
	CUT_1711:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(11));
	CUT_1712:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(12));
	CUT_1713:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(13));
	CUT_1714:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(14));
	CUT_1715:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(15));
	CUT_1716:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(16));
	CUT_1717:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(17));
	CUT_1718:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(18));
	CUT_1719:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(19));
	CUT_1720:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(20));
	CUT_1721:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(21));
	CUT_1722:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(22));
	CUT_1723:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(23));
	CUT_1724:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(24));
	CUT_1725:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(25));
	CUT_1726:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(26));
	CUT_1727:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(27));
	CUT_1728:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(28));
	CUT_1729:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(29));
	CUT_1730:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(30));
	CUT_1731:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(31));
	CUT_1732:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(32));
	CUT_1733:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(33));
	CUT_1734:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(34));
	CUT_1735:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(35));
	CUT_1736:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(36));
	CUT_1737:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(37));
	CUT_1738:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(38));
	CUT_1739:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(39));
	CUT_1740:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(40));
	CUT_1741:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(41));
	CUT_1742:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(42));
	CUT_1743:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(43));
	CUT_1744:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(44));
	CUT_1745:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(45));
	CUT_1746:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(46));
	CUT_1747:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(47));
	CUT_1748:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(48));
	CUT_1749:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(34)(49));
	CUT_1750:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(0));
	CUT_1751:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(1));
	CUT_1752:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(2));
	CUT_1753:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(3));
	CUT_1754:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(4));
	CUT_1755:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(5));
	CUT_1756:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(6));
	CUT_1757:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(7));
	CUT_1758:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(8));
	CUT_1759:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(9));
	CUT_1760:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(10));
	CUT_1761:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(11));
	CUT_1762:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(12));
	CUT_1763:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(13));
	CUT_1764:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(14));
	CUT_1765:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(15));
	CUT_1766:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(16));
	CUT_1767:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(17));
	CUT_1768:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(18));
	CUT_1769:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(19));
	CUT_1770:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(20));
	CUT_1771:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(21));
	CUT_1772:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(22));
	CUT_1773:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(23));
	CUT_1774:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(24));
	CUT_1775:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(25));
	CUT_1776:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(26));
	CUT_1777:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(27));
	CUT_1778:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(28));
	CUT_1779:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(29));
	CUT_1780:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(30));
	CUT_1781:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(31));
	CUT_1782:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(32));
	CUT_1783:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(33));
	CUT_1784:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(34));
	CUT_1785:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(35));
	CUT_1786:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(36));
	CUT_1787:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(37));
	CUT_1788:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(38));
	CUT_1789:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(39));
	CUT_1790:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(40));
	CUT_1791:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(41));
	CUT_1792:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(42));
	CUT_1793:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(43));
	CUT_1794:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(44));
	CUT_1795:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(45));
	CUT_1796:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(46));
	CUT_1797:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(47));
	CUT_1798:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(48));
	CUT_1799:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(35)(49));
	CUT_1800:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(0));
	CUT_1801:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(1));
	CUT_1802:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(2));
	CUT_1803:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(3));
	CUT_1804:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(4));
	CUT_1805:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(5));
	CUT_1806:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(6));
	CUT_1807:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(7));
	CUT_1808:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(8));
	CUT_1809:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(9));
	CUT_1810:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(10));
	CUT_1811:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(11));
	CUT_1812:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(12));
	CUT_1813:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(13));
	CUT_1814:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(14));
	CUT_1815:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(15));
	CUT_1816:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(16));
	CUT_1817:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(17));
	CUT_1818:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(18));
	CUT_1819:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(19));
	CUT_1820:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(20));
	CUT_1821:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(21));
	CUT_1822:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(22));
	CUT_1823:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(23));
	CUT_1824:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(24));
	CUT_1825:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(25));
	CUT_1826:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(26));
	CUT_1827:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(27));
	CUT_1828:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(28));
	CUT_1829:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(29));
	CUT_1830:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(30));
	CUT_1831:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(31));
	CUT_1832:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(32));
	CUT_1833:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(33));
	CUT_1834:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(34));
	CUT_1835:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(35));
	CUT_1836:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(36));
	CUT_1837:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(37));
	CUT_1838:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(38));
	CUT_1839:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(39));
	CUT_1840:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(40));
	CUT_1841:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(41));
	CUT_1842:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(42));
	CUT_1843:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(43));
	CUT_1844:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(44));
	CUT_1845:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(45));
	CUT_1846:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(46));
	CUT_1847:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(47));
	CUT_1848:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(48));
	CUT_1849:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(36)(49));
	CUT_1850:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(0));
	CUT_1851:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(1));
	CUT_1852:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(2));
	CUT_1853:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(3));
	CUT_1854:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(4));
	CUT_1855:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(5));
	CUT_1856:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(6));
	CUT_1857:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(7));
	CUT_1858:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(8));
	CUT_1859:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(9));
	CUT_1860:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(10));
	CUT_1861:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(11));
	CUT_1862:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(12));
	CUT_1863:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(13));
	CUT_1864:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(14));
	CUT_1865:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(15));
	CUT_1866:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(16));
	CUT_1867:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(17));
	CUT_1868:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(18));
	CUT_1869:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(19));
	CUT_1870:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(20));
	CUT_1871:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(21));
	CUT_1872:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(22));
	CUT_1873:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(23));
	CUT_1874:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(24));
	CUT_1875:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(25));
	CUT_1876:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(26));
	CUT_1877:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(27));
	CUT_1878:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(28));
	CUT_1879:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(29));
	CUT_1880:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(30));
	CUT_1881:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(31));
	CUT_1882:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(32));
	CUT_1883:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(33));
	CUT_1884:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(34));
	CUT_1885:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(35));
	CUT_1886:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(36));
	CUT_1887:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(37));
	CUT_1888:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(38));
	CUT_1889:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(39));
	CUT_1890:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(40));
	CUT_1891:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(41));
	CUT_1892:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(42));
	CUT_1893:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(43));
	CUT_1894:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(44));
	CUT_1895:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(45));
	CUT_1896:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(46));
	CUT_1897:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(47));
	CUT_1898:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(48));
	CUT_1899:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(37)(49));
	CUT_1900:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(0));
	CUT_1901:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(1));
	CUT_1902:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(2));
	CUT_1903:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(3));
	CUT_1904:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(4));
	CUT_1905:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(5));
	CUT_1906:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(6));
	CUT_1907:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(7));
	CUT_1908:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(8));
	CUT_1909:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(9));
	CUT_1910:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(10));
	CUT_1911:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(11));
	CUT_1912:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(12));
	CUT_1913:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(13));
	CUT_1914:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(14));
	CUT_1915:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(15));
	CUT_1916:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(16));
	CUT_1917:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(17));
	CUT_1918:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(18));
	CUT_1919:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(19));
	CUT_1920:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(20));
	CUT_1921:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(21));
	CUT_1922:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(22));
	CUT_1923:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(23));
	CUT_1924:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(24));
	CUT_1925:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(25));
	CUT_1926:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(26));
	CUT_1927:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(27));
	CUT_1928:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(28));
	CUT_1929:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(29));
	CUT_1930:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(30));
	CUT_1931:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(31));
	CUT_1932:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(32));
	CUT_1933:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(33));
	CUT_1934:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(34));
	CUT_1935:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(35));
	CUT_1936:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(36));
	CUT_1937:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(37));
	CUT_1938:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(38));
	CUT_1939:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(39));
	CUT_1940:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(40));
	CUT_1941:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(41));
	CUT_1942:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(42));
	CUT_1943:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(43));
	CUT_1944:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(44));
	CUT_1945:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(45));
	CUT_1946:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(46));
	CUT_1947:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(47));
	CUT_1948:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(48));
	CUT_1949:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(38)(49));
	CUT_1950:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(0));
	CUT_1951:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(1));
	CUT_1952:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(2));
	CUT_1953:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(3));
	CUT_1954:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(4));
	CUT_1955:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(5));
	CUT_1956:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(6));
	CUT_1957:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(7));
	CUT_1958:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(8));
	CUT_1959:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(9));
	CUT_1960:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(10));
	CUT_1961:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(11));
	CUT_1962:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(12));
	CUT_1963:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(13));
	CUT_1964:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(14));
	CUT_1965:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(15));
	CUT_1966:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(16));
	CUT_1967:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(17));
	CUT_1968:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(18));
	CUT_1969:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(19));
	CUT_1970:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(20));
	CUT_1971:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(21));
	CUT_1972:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(22));
	CUT_1973:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(23));
	CUT_1974:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(24));
	CUT_1975:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(25));
	CUT_1976:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(26));
	CUT_1977:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(27));
	CUT_1978:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(28));
	CUT_1979:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(29));
	CUT_1980:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(30));
	CUT_1981:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(31));
	CUT_1982:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(32));
	CUT_1983:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(33));
	CUT_1984:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(34));
	CUT_1985:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(35));
	CUT_1986:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(36));
	CUT_1987:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(37));
	CUT_1988:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(38));
	CUT_1989:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(39));
	CUT_1990:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(40));
	CUT_1991:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(41));
	CUT_1992:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(42));
	CUT_1993:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(43));
	CUT_1994:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(44));
	CUT_1995:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(45));
	CUT_1996:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(46));
	CUT_1997:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(47));
	CUT_1998:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(48));
	CUT_1999:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(39)(49));
	CUT_2000:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(0));
	CUT_2001:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(1));
	CUT_2002:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(2));
	CUT_2003:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(3));
	CUT_2004:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(4));
	CUT_2005:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(5));
	CUT_2006:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(6));
	CUT_2007:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(7));
	CUT_2008:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(8));
	CUT_2009:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(9));
	CUT_2010:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(10));
	CUT_2011:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(11));
	CUT_2012:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(12));
	CUT_2013:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(13));
	CUT_2014:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(14));
	CUT_2015:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(15));
	CUT_2016:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(16));
	CUT_2017:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(17));
	CUT_2018:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(18));
	CUT_2019:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(19));
	CUT_2020:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(20));
	CUT_2021:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(21));
	CUT_2022:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(22));
	CUT_2023:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(23));
	CUT_2024:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(24));
	CUT_2025:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(25));
	CUT_2026:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(26));
	CUT_2027:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(27));
	CUT_2028:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(28));
	CUT_2029:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(29));
	CUT_2030:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(30));
	CUT_2031:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(31));
	CUT_2032:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(32));
	CUT_2033:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(33));
	CUT_2034:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(34));
	CUT_2035:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(35));
	CUT_2036:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(36));
	CUT_2037:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(37));
	CUT_2038:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(38));
	CUT_2039:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(39));
	CUT_2040:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(40));
	CUT_2041:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(41));
	CUT_2042:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(42));
	CUT_2043:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(43));
	CUT_2044:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(44));
	CUT_2045:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(45));
	CUT_2046:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(46));
	CUT_2047:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(47));
	CUT_2048:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(48));
	CUT_2049:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(40)(49));
	CUT_2050:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(0));
	CUT_2051:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(1));
	CUT_2052:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(2));
	CUT_2053:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(3));
	CUT_2054:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(4));
	CUT_2055:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(5));
	CUT_2056:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(6));
	CUT_2057:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(7));
	CUT_2058:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(8));
	CUT_2059:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(9));
	CUT_2060:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(10));
	CUT_2061:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(11));
	CUT_2062:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(12));
	CUT_2063:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(13));
	CUT_2064:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(14));
	CUT_2065:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(15));
	CUT_2066:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(16));
	CUT_2067:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(17));
	CUT_2068:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(18));
	CUT_2069:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(19));
	CUT_2070:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(20));
	CUT_2071:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(21));
	CUT_2072:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(22));
	CUT_2073:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(23));
	CUT_2074:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(24));
	CUT_2075:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(25));
	CUT_2076:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(26));
	CUT_2077:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(27));
	CUT_2078:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(28));
	CUT_2079:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(29));
	CUT_2080:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(30));
	CUT_2081:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(31));
	CUT_2082:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(32));
	CUT_2083:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(33));
	CUT_2084:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(34));
	CUT_2085:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(35));
	CUT_2086:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(36));
	CUT_2087:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(37));
	CUT_2088:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(38));
	CUT_2089:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(39));
	CUT_2090:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(40));
	CUT_2091:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(41));
	CUT_2092:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(42));
	CUT_2093:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(43));
	CUT_2094:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(44));
	CUT_2095:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(45));
	CUT_2096:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(46));
	CUT_2097:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(47));
	CUT_2098:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(48));
	CUT_2099:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(41)(49));
	CUT_2100:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(0));
	CUT_2101:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(1));
	CUT_2102:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(2));
	CUT_2103:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(3));
	CUT_2104:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(4));
	CUT_2105:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(5));
	CUT_2106:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(6));
	CUT_2107:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(7));
	CUT_2108:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(8));
	CUT_2109:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(9));
	CUT_2110:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(10));
	CUT_2111:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(11));
	CUT_2112:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(12));
	CUT_2113:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(13));
	CUT_2114:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(14));
	CUT_2115:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(15));
	CUT_2116:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(16));
	CUT_2117:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(17));
	CUT_2118:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(18));
	CUT_2119:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(19));
	CUT_2120:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(20));
	CUT_2121:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(21));
	CUT_2122:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(22));
	CUT_2123:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(23));
	CUT_2124:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(24));
	CUT_2125:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(25));
	CUT_2126:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(26));
	CUT_2127:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(27));
	CUT_2128:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(28));
	CUT_2129:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(29));
	CUT_2130:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(30));
	CUT_2131:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(31));
	CUT_2132:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(32));
	CUT_2133:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(33));
	CUT_2134:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(34));
	CUT_2135:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(35));
	CUT_2136:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(36));
	CUT_2137:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(37));
	CUT_2138:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(38));
	CUT_2139:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(39));
	CUT_2140:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(40));
	CUT_2141:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(41));
	CUT_2142:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(42));
	CUT_2143:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(43));
	CUT_2144:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(44));
	CUT_2145:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(45));
	CUT_2146:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(46));
	CUT_2147:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(47));
	CUT_2148:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(48));
	CUT_2149:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(42)(49));
	CUT_2150:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(0));
	CUT_2151:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(1));
	CUT_2152:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(2));
	CUT_2153:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(3));
	CUT_2154:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(4));
	CUT_2155:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(5));
	CUT_2156:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(6));
	CUT_2157:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(7));
	CUT_2158:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(8));
	CUT_2159:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(9));
	CUT_2160:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(10));
	CUT_2161:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(11));
	CUT_2162:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(12));
	CUT_2163:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(13));
	CUT_2164:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(14));
	CUT_2165:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(15));
	CUT_2166:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(16));
	CUT_2167:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(17));
	CUT_2168:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(18));
	CUT_2169:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(19));
	CUT_2170:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(20));
	CUT_2171:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(21));
	CUT_2172:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(22));
	CUT_2173:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(23));
	CUT_2174:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(24));
	CUT_2175:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(25));
	CUT_2176:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(26));
	CUT_2177:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(27));
	CUT_2178:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(28));
	CUT_2179:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(29));
	CUT_2180:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(30));
	CUT_2181:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(31));
	CUT_2182:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(32));
	CUT_2183:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(33));
	CUT_2184:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(34));
	CUT_2185:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(35));
	CUT_2186:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(36));
	CUT_2187:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(37));
	CUT_2188:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(38));
	CUT_2189:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(39));
	CUT_2190:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(40));
	CUT_2191:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(41));
	CUT_2192:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(42));
	CUT_2193:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(43));
	CUT_2194:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(44));
	CUT_2195:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(45));
	CUT_2196:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(46));
	CUT_2197:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(47));
	CUT_2198:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(48));
	CUT_2199:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(43)(49));
	CUT_2200:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(0));
	CUT_2201:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(1));
	CUT_2202:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(2));
	CUT_2203:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(3));
	CUT_2204:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(4));
	CUT_2205:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(5));
	CUT_2206:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(6));
	CUT_2207:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(7));
	CUT_2208:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(8));
	CUT_2209:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(9));
	CUT_2210:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(10));
	CUT_2211:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(11));
	CUT_2212:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(12));
	CUT_2213:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(13));
	CUT_2214:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(14));
	CUT_2215:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(15));
	CUT_2216:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(16));
	CUT_2217:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(17));
	CUT_2218:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(18));
	CUT_2219:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(19));
	CUT_2220:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(20));
	CUT_2221:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(21));
	CUT_2222:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(22));
	CUT_2223:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(23));
	CUT_2224:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(24));
	CUT_2225:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(25));
	CUT_2226:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(26));
	CUT_2227:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(27));
	CUT_2228:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(28));
	CUT_2229:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(29));
	CUT_2230:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(30));
	CUT_2231:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(31));
	CUT_2232:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(32));
	CUT_2233:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(33));
	CUT_2234:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(34));
	CUT_2235:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(35));
	CUT_2236:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(36));
	CUT_2237:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(37));
	CUT_2238:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(38));
	CUT_2239:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(39));
	CUT_2240:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(40));
	CUT_2241:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(41));
	CUT_2242:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(42));
	CUT_2243:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(43));
	CUT_2244:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(44));
	CUT_2245:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(45));
	CUT_2246:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(46));
	CUT_2247:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(47));
	CUT_2248:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(48));
	CUT_2249:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(44)(49));
	CUT_2250:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(0));
	CUT_2251:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(1));
	CUT_2252:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(2));
	CUT_2253:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(3));
	CUT_2254:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(4));
	CUT_2255:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(5));
	CUT_2256:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(6));
	CUT_2257:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(7));
	CUT_2258:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(8));
	CUT_2259:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(9));
	CUT_2260:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(10));
	CUT_2261:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(11));
	CUT_2262:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(12));
	CUT_2263:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(13));
	CUT_2264:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(14));
	CUT_2265:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(15));
	CUT_2266:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(16));
	CUT_2267:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(17));
	CUT_2268:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(18));
	CUT_2269:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(19));
	CUT_2270:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(20));
	CUT_2271:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(21));
	CUT_2272:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(22));
	CUT_2273:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(23));
	CUT_2274:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(24));
	CUT_2275:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(25));
	CUT_2276:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(26));
	CUT_2277:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(27));
	CUT_2278:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(28));
	CUT_2279:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(29));
	CUT_2280:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(30));
	CUT_2281:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(31));
	CUT_2282:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(32));
	CUT_2283:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(33));
	CUT_2284:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(34));
	CUT_2285:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(35));
	CUT_2286:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(36));
	CUT_2287:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(37));
	CUT_2288:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(38));
	CUT_2289:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(39));
	CUT_2290:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(40));
	CUT_2291:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(41));
	CUT_2292:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(42));
	CUT_2293:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(43));
	CUT_2294:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(44));
	CUT_2295:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(45));
	CUT_2296:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(46));
	CUT_2297:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(47));
	CUT_2298:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(48));
	CUT_2299:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(45)(49));
	CUT_2300:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(0));
	CUT_2301:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(1));
	CUT_2302:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(2));
	CUT_2303:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(3));
	CUT_2304:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(4));
	CUT_2305:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(5));
	CUT_2306:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(6));
	CUT_2307:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(7));
	CUT_2308:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(8));
	CUT_2309:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(9));
	CUT_2310:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(10));
	CUT_2311:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(11));
	CUT_2312:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(12));
	CUT_2313:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(13));
	CUT_2314:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(14));
	CUT_2315:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(15));
	CUT_2316:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(16));
	CUT_2317:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(17));
	CUT_2318:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(18));
	CUT_2319:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(19));
	CUT_2320:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(20));
	CUT_2321:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(21));
	CUT_2322:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(22));
	CUT_2323:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(23));
	CUT_2324:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(24));
	CUT_2325:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(25));
	CUT_2326:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(26));
	CUT_2327:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(27));
	CUT_2328:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(28));
	CUT_2329:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(29));
	CUT_2330:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(30));
	CUT_2331:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(31));
	CUT_2332:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(32));
	CUT_2333:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(33));
	CUT_2334:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(34));
	CUT_2335:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(35));
	CUT_2336:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(36));
	CUT_2337:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(37));
	CUT_2338:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(38));
	CUT_2339:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(39));
	CUT_2340:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(40));
	CUT_2341:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(41));
	CUT_2342:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(42));
	CUT_2343:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(43));
	CUT_2344:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(44));
	CUT_2345:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(45));
	CUT_2346:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(46));
	CUT_2347:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(47));
	CUT_2348:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(48));
	CUT_2349:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(46)(49));
	CUT_2350:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(0));
	CUT_2351:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(1));
	CUT_2352:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(2));
	CUT_2353:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(3));
	CUT_2354:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(4));
	CUT_2355:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(5));
	CUT_2356:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(6));
	CUT_2357:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(7));
	CUT_2358:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(8));
	CUT_2359:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(9));
	CUT_2360:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(10));
	CUT_2361:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(11));
	CUT_2362:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(12));
	CUT_2363:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(13));
	CUT_2364:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(14));
	CUT_2365:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(15));
	CUT_2366:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(16));
	CUT_2367:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(17));
	CUT_2368:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(18));
	CUT_2369:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(19));
	CUT_2370:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(20));
	CUT_2371:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(21));
	CUT_2372:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(22));
	CUT_2373:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(23));
	CUT_2374:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(24));
	CUT_2375:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(25));
	CUT_2376:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(26));
	CUT_2377:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(27));
	CUT_2378:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(28));
	CUT_2379:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(29));
	CUT_2380:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(30));
	CUT_2381:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(31));
	CUT_2382:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(32));
	CUT_2383:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(33));
	CUT_2384:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(34));
	CUT_2385:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(35));
	CUT_2386:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(36));
	CUT_2387:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(37));
	CUT_2388:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(38));
	CUT_2389:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(39));
	CUT_2390:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(40));
	CUT_2391:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(41));
	CUT_2392:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(42));
	CUT_2393:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(43));
	CUT_2394:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(44));
	CUT_2395:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(45));
	CUT_2396:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(46));
	CUT_2397:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(47));
	CUT_2398:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(48));
	CUT_2399:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(47)(49));
	CUT_2400:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(0));
	CUT_2401:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(1));
	CUT_2402:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(2));
	CUT_2403:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(3));
	CUT_2404:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(4));
	CUT_2405:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(5));
	CUT_2406:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(6));
	CUT_2407:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(7));
	CUT_2408:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(8));
	CUT_2409:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(9));
	CUT_2410:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(10));
	CUT_2411:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(11));
	CUT_2412:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(12));
	CUT_2413:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(13));
	CUT_2414:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(14));
	CUT_2415:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(15));
	CUT_2416:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(16));
	CUT_2417:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(17));
	CUT_2418:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(18));
	CUT_2419:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(19));
	CUT_2420:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(20));
	CUT_2421:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(21));
	CUT_2422:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(22));
	CUT_2423:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(23));
	CUT_2424:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(24));
	CUT_2425:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(25));
	CUT_2426:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(26));
	CUT_2427:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(27));
	CUT_2428:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(28));
	CUT_2429:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(29));
	CUT_2430:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(30));
	CUT_2431:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(31));
	CUT_2432:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(32));
	CUT_2433:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(33));
	CUT_2434:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(34));
	CUT_2435:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(35));
	CUT_2436:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(36));
	CUT_2437:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(37));
	CUT_2438:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(38));
	CUT_2439:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(39));
	CUT_2440:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(40));
	CUT_2441:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(41));
	CUT_2442:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(42));
	CUT_2443:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(43));
	CUT_2444:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(44));
	CUT_2445:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(45));
	CUT_2446:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(46));
	CUT_2447:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(47));
	CUT_2448:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(48));
	CUT_2449:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(48)(49));
	CUT_2450:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(0));
	CUT_2451:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(1));
	CUT_2452:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(2));
	CUT_2453:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(3));
	CUT_2454:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(4));
	CUT_2455:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(5));
	CUT_2456:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(6));
	CUT_2457:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(7));
	CUT_2458:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(8));
	CUT_2459:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(9));
	CUT_2460:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(10));
	CUT_2461:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(11));
	CUT_2462:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(12));
	CUT_2463:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(13));
	CUT_2464:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(14));
	CUT_2465:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(15));
	CUT_2466:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(16));
	CUT_2467:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(17));
	CUT_2468:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(18));
	CUT_2469:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(19));
	CUT_2470:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(20));
	CUT_2471:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(21));
	CUT_2472:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(22));
	CUT_2473:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(23));
	CUT_2474:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(24));
	CUT_2475:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(25));
	CUT_2476:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(26));
	CUT_2477:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(27));
	CUT_2478:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(28));
	CUT_2479:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(29));
	CUT_2480:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(30));
	CUT_2481:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(31));
	CUT_2482:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(32));
	CUT_2483:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(33));
	CUT_2484:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(34));
	CUT_2485:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(35));
	CUT_2486:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(36));
	CUT_2487:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(37));
	CUT_2488:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(38));
	CUT_2489:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(39));
	CUT_2490:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(40));
	CUT_2491:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(41));
	CUT_2492:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(42));
	CUT_2493:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(43));
	CUT_2494:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(44));
	CUT_2495:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(45));
	CUT_2496:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(46));
	CUT_2497:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(47));
	CUT_2498:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(48));
	CUT_2499:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(49)(49));
	CUT_2500:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(0));
	CUT_2501:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(1));
	CUT_2502:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(2));
	CUT_2503:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(3));
	CUT_2504:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(4));
	CUT_2505:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(5));
	CUT_2506:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(6));
	CUT_2507:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(7));
	CUT_2508:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(8));
	CUT_2509:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(9));
	CUT_2510:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(10));
	CUT_2511:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(11));
	CUT_2512:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(12));
	CUT_2513:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(13));
	CUT_2514:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(14));
	CUT_2515:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(15));
	CUT_2516:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(16));
	CUT_2517:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(17));
	CUT_2518:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(18));
	CUT_2519:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(19));
	CUT_2520:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(20));
	CUT_2521:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(21));
	CUT_2522:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(22));
	CUT_2523:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(23));
	CUT_2524:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(24));
	CUT_2525:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(25));
	CUT_2526:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(26));
	CUT_2527:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(27));
	CUT_2528:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(28));
	CUT_2529:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(29));
	CUT_2530:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(30));
	CUT_2531:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(31));
	CUT_2532:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(32));
	CUT_2533:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(33));
	CUT_2534:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(34));
	CUT_2535:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(35));
	CUT_2536:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(36));
	CUT_2537:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(37));
	CUT_2538:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(38));
	CUT_2539:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(39));
	CUT_2540:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(40));
	CUT_2541:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(41));
	CUT_2542:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(42));
	CUT_2543:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(43));
	CUT_2544:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(44));
	CUT_2545:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(45));
	CUT_2546:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(46));
	CUT_2547:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(47));
	CUT_2548:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(48));
	CUT_2549:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(50)(49));
	CUT_2550:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(0));
	CUT_2551:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(1));
	CUT_2552:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(2));
	CUT_2553:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(3));
	CUT_2554:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(4));
	CUT_2555:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(5));
	CUT_2556:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(6));
	CUT_2557:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(7));
	CUT_2558:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(8));
	CUT_2559:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(9));
	CUT_2560:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(10));
	CUT_2561:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(11));
	CUT_2562:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(12));
	CUT_2563:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(13));
	CUT_2564:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(14));
	CUT_2565:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(15));
	CUT_2566:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(16));
	CUT_2567:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(17));
	CUT_2568:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(18));
	CUT_2569:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(19));
	CUT_2570:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(20));
	CUT_2571:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(21));
	CUT_2572:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(22));
	CUT_2573:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(23));
	CUT_2574:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(24));
	CUT_2575:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(25));
	CUT_2576:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(26));
	CUT_2577:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(27));
	CUT_2578:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(28));
	CUT_2579:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(29));
	CUT_2580:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(30));
	CUT_2581:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(31));
	CUT_2582:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(32));
	CUT_2583:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(33));
	CUT_2584:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(34));
	CUT_2585:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(35));
	CUT_2586:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(36));
	CUT_2587:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(37));
	CUT_2588:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(38));
	CUT_2589:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(39));
	CUT_2590:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(40));
	CUT_2591:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(41));
	CUT_2592:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(42));
	CUT_2593:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(43));
	CUT_2594:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(44));
	CUT_2595:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(45));
	CUT_2596:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(46));
	CUT_2597:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(47));
	CUT_2598:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(48));
	CUT_2599:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(51)(49));
	CUT_2600:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(0));
	CUT_2601:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(1));
	CUT_2602:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(2));
	CUT_2603:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(3));
	CUT_2604:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(4));
	CUT_2605:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(5));
	CUT_2606:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(6));
	CUT_2607:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(7));
	CUT_2608:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(8));
	CUT_2609:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(9));
	CUT_2610:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(10));
	CUT_2611:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(11));
	CUT_2612:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(12));
	CUT_2613:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(13));
	CUT_2614:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(14));
	CUT_2615:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(15));
	CUT_2616:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(16));
	CUT_2617:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(17));
	CUT_2618:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(18));
	CUT_2619:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(19));
	CUT_2620:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(20));
	CUT_2621:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(21));
	CUT_2622:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(22));
	CUT_2623:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(23));
	CUT_2624:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(24));
	CUT_2625:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(25));
	CUT_2626:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(26));
	CUT_2627:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(27));
	CUT_2628:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(28));
	CUT_2629:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(29));
	CUT_2630:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(30));
	CUT_2631:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(31));
	CUT_2632:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(32));
	CUT_2633:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(33));
	CUT_2634:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(34));
	CUT_2635:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(35));
	CUT_2636:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(36));
	CUT_2637:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(37));
	CUT_2638:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(38));
	CUT_2639:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(39));
	CUT_2640:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(40));
	CUT_2641:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(41));
	CUT_2642:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(42));
	CUT_2643:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(43));
	CUT_2644:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(44));
	CUT_2645:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(45));
	CUT_2646:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(46));
	CUT_2647:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(47));
	CUT_2648:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(48));
	CUT_2649:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(52)(49));
	CUT_2650:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(0));
	CUT_2651:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(1));
	CUT_2652:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(2));
	CUT_2653:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(3));
	CUT_2654:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(4));
	CUT_2655:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(5));
	CUT_2656:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(6));
	CUT_2657:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(7));
	CUT_2658:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(8));
	CUT_2659:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(9));
	CUT_2660:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(10));
	CUT_2661:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(11));
	CUT_2662:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(12));
	CUT_2663:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(13));
	CUT_2664:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(14));
	CUT_2665:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(15));
	CUT_2666:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(16));
	CUT_2667:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(17));
	CUT_2668:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(18));
	CUT_2669:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(19));
	CUT_2670:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(20));
	CUT_2671:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(21));
	CUT_2672:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(22));
	CUT_2673:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(23));
	CUT_2674:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(24));
	CUT_2675:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(25));
	CUT_2676:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(26));
	CUT_2677:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(27));
	CUT_2678:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(28));
	CUT_2679:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(29));
	CUT_2680:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(30));
	CUT_2681:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(31));
	CUT_2682:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(32));
	CUT_2683:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(33));
	CUT_2684:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(34));
	CUT_2685:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(35));
	CUT_2686:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(36));
	CUT_2687:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(37));
	CUT_2688:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(38));
	CUT_2689:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(39));
	CUT_2690:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(40));
	CUT_2691:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(41));
	CUT_2692:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(42));
	CUT_2693:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(43));
	CUT_2694:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(44));
	CUT_2695:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(45));
	CUT_2696:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(46));
	CUT_2697:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(47));
	CUT_2698:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(48));
	CUT_2699:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(53)(49));
	CUT_2700:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(0));
	CUT_2701:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(1));
	CUT_2702:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(2));
	CUT_2703:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(3));
	CUT_2704:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(4));
	CUT_2705:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(5));
	CUT_2706:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(6));
	CUT_2707:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(7));
	CUT_2708:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(8));
	CUT_2709:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(9));
	CUT_2710:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(10));
	CUT_2711:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(11));
	CUT_2712:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(12));
	CUT_2713:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(13));
	CUT_2714:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(14));
	CUT_2715:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(15));
	CUT_2716:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(16));
	CUT_2717:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(17));
	CUT_2718:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(18));
	CUT_2719:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(19));
	CUT_2720:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(20));
	CUT_2721:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(21));
	CUT_2722:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(22));
	CUT_2723:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(23));
	CUT_2724:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(24));
	CUT_2725:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(25));
	CUT_2726:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(26));
	CUT_2727:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(27));
	CUT_2728:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(28));
	CUT_2729:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(29));
	CUT_2730:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(30));
	CUT_2731:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(31));
	CUT_2732:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(32));
	CUT_2733:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(33));
	CUT_2734:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(34));
	CUT_2735:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(35));
	CUT_2736:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(36));
	CUT_2737:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(37));
	CUT_2738:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(38));
	CUT_2739:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(39));
	CUT_2740:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(40));
	CUT_2741:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(41));
	CUT_2742:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(42));
	CUT_2743:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(43));
	CUT_2744:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(44));
	CUT_2745:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(45));
	CUT_2746:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(46));
	CUT_2747:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(47));
	CUT_2748:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(48));
	CUT_2749:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(54)(49));
	CUT_2750:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(0));
	CUT_2751:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(1));
	CUT_2752:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(2));
	CUT_2753:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(3));
	CUT_2754:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(4));
	CUT_2755:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(5));
	CUT_2756:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(6));
	CUT_2757:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(7));
	CUT_2758:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(8));
	CUT_2759:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(9));
	CUT_2760:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(10));
	CUT_2761:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(11));
	CUT_2762:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(12));
	CUT_2763:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(13));
	CUT_2764:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(14));
	CUT_2765:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(15));
	CUT_2766:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(16));
	CUT_2767:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(17));
	CUT_2768:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(18));
	CUT_2769:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(19));
	CUT_2770:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(20));
	CUT_2771:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(21));
	CUT_2772:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(22));
	CUT_2773:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(23));
	CUT_2774:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(24));
	CUT_2775:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(25));
	CUT_2776:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(26));
	CUT_2777:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(27));
	CUT_2778:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(28));
	CUT_2779:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(29));
	CUT_2780:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(30));
	CUT_2781:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(31));
	CUT_2782:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(32));
	CUT_2783:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(33));
	CUT_2784:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(34));
	CUT_2785:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(35));
	CUT_2786:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(36));
	CUT_2787:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(37));
	CUT_2788:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(38));
	CUT_2789:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(39));
	CUT_2790:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(40));
	CUT_2791:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(41));
	CUT_2792:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(42));
	CUT_2793:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(43));
	CUT_2794:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(44));
	CUT_2795:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(45));
	CUT_2796:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(46));
	CUT_2797:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(47));
	CUT_2798:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(48));
	CUT_2799:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(55)(49));
	CUT_2800:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(0));
	CUT_2801:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(1));
	CUT_2802:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(2));
	CUT_2803:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(3));
	CUT_2804:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(4));
	CUT_2805:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(5));
	CUT_2806:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(6));
	CUT_2807:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(7));
	CUT_2808:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(8));
	CUT_2809:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(9));
	CUT_2810:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(10));
	CUT_2811:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(11));
	CUT_2812:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(12));
	CUT_2813:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(13));
	CUT_2814:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(14));
	CUT_2815:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(15));
	CUT_2816:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(16));
	CUT_2817:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(17));
	CUT_2818:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(18));
	CUT_2819:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(19));
	CUT_2820:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(20));
	CUT_2821:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(21));
	CUT_2822:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(22));
	CUT_2823:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(23));
	CUT_2824:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(24));
	CUT_2825:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(25));
	CUT_2826:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(26));
	CUT_2827:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(27));
	CUT_2828:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(28));
	CUT_2829:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(29));
	CUT_2830:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(30));
	CUT_2831:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(31));
	CUT_2832:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(32));
	CUT_2833:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(33));
	CUT_2834:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(34));
	CUT_2835:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(35));
	CUT_2836:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(36));
	CUT_2837:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(37));
	CUT_2838:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(38));
	CUT_2839:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(39));
	CUT_2840:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(40));
	CUT_2841:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(41));
	CUT_2842:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(42));
	CUT_2843:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(43));
	CUT_2844:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(44));
	CUT_2845:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(45));
	CUT_2846:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(46));
	CUT_2847:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(47));
	CUT_2848:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(48));
	CUT_2849:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(56)(49));
	CUT_2850:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(0));
	CUT_2851:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(1));
	CUT_2852:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(2));
	CUT_2853:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(3));
	CUT_2854:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(4));
	CUT_2855:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(5));
	CUT_2856:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(6));
	CUT_2857:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(7));
	CUT_2858:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(8));
	CUT_2859:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(9));
	CUT_2860:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(10));
	CUT_2861:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(11));
	CUT_2862:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(12));
	CUT_2863:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(13));
	CUT_2864:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(14));
	CUT_2865:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(15));
	CUT_2866:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(16));
	CUT_2867:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(17));
	CUT_2868:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(18));
	CUT_2869:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(19));
	CUT_2870:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(20));
	CUT_2871:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(21));
	CUT_2872:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(22));
	CUT_2873:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(23));
	CUT_2874:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(24));
	CUT_2875:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(25));
	CUT_2876:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(26));
	CUT_2877:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(27));
	CUT_2878:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(28));
	CUT_2879:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(29));
	CUT_2880:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(30));
	CUT_2881:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(31));
	CUT_2882:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(32));
	CUT_2883:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(33));
	CUT_2884:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(34));
	CUT_2885:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(35));
	CUT_2886:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(36));
	CUT_2887:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(37));
	CUT_2888:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(38));
	CUT_2889:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(39));
	CUT_2890:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(40));
	CUT_2891:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(41));
	CUT_2892:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(42));
	CUT_2893:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(43));
	CUT_2894:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(44));
	CUT_2895:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(45));
	CUT_2896:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(46));
	CUT_2897:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(47));
	CUT_2898:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(48));
	CUT_2899:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(57)(49));
	CUT_2900:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(0));
	CUT_2901:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(1));
	CUT_2902:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(2));
	CUT_2903:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(3));
	CUT_2904:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(4));
	CUT_2905:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(5));
	CUT_2906:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(6));
	CUT_2907:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(7));
	CUT_2908:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(8));
	CUT_2909:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(9));
	CUT_2910:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(10));
	CUT_2911:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(11));
	CUT_2912:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(12));
	CUT_2913:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(13));
	CUT_2914:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(14));
	CUT_2915:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(15));
	CUT_2916:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(16));
	CUT_2917:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(17));
	CUT_2918:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(18));
	CUT_2919:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(19));
	CUT_2920:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(20));
	CUT_2921:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(21));
	CUT_2922:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(22));
	CUT_2923:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(23));
	CUT_2924:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(24));
	CUT_2925:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(25));
	CUT_2926:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(26));
	CUT_2927:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(27));
	CUT_2928:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(28));
	CUT_2929:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(29));
	CUT_2930:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(30));
	CUT_2931:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(31));
	CUT_2932:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(32));
	CUT_2933:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(33));
	CUT_2934:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(34));
	CUT_2935:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(35));
	CUT_2936:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(36));
	CUT_2937:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(37));
	CUT_2938:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(38));
	CUT_2939:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(39));
	CUT_2940:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(40));
	CUT_2941:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(41));
	CUT_2942:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(42));
	CUT_2943:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(43));
	CUT_2944:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(44));
	CUT_2945:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(45));
	CUT_2946:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(46));
	CUT_2947:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(47));
	CUT_2948:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(48));
	CUT_2949:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(58)(49));
	CUT_2950:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(0));
	CUT_2951:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(1));
	CUT_2952:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(2));
	CUT_2953:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(3));
	CUT_2954:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(4));
	CUT_2955:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(5));
	CUT_2956:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(6));
	CUT_2957:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(7));
	CUT_2958:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(8));
	CUT_2959:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(9));
	CUT_2960:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(10));
	CUT_2961:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(11));
	CUT_2962:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(12));
	CUT_2963:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(13));
	CUT_2964:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(14));
	CUT_2965:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(15));
	CUT_2966:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(16));
	CUT_2967:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(17));
	CUT_2968:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(18));
	CUT_2969:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(19));
	CUT_2970:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(20));
	CUT_2971:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(21));
	CUT_2972:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(22));
	CUT_2973:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(23));
	CUT_2974:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(24));
	CUT_2975:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(25));
	CUT_2976:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(26));
	CUT_2977:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(27));
	CUT_2978:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(28));
	CUT_2979:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(29));
	CUT_2980:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(30));
	CUT_2981:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(31));
	CUT_2982:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(32));
	CUT_2983:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(33));
	CUT_2984:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(34));
	CUT_2985:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(35));
	CUT_2986:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(36));
	CUT_2987:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(37));
	CUT_2988:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(38));
	CUT_2989:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(39));
	CUT_2990:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(40));
	CUT_2991:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(41));
	CUT_2992:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(42));
	CUT_2993:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(43));
	CUT_2994:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(44));
	CUT_2995:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(45));
	CUT_2996:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(46));
	CUT_2997:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(47));
	CUT_2998:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(48));
	CUT_2999:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(59)(49));
	CUT_3000:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(0));
	CUT_3001:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(1));
	CUT_3002:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(2));
	CUT_3003:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(3));
	CUT_3004:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(4));
	CUT_3005:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(5));
	CUT_3006:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(6));
	CUT_3007:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(7));
	CUT_3008:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(8));
	CUT_3009:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(9));
	CUT_3010:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(10));
	CUT_3011:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(11));
	CUT_3012:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(12));
	CUT_3013:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(13));
	CUT_3014:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(14));
	CUT_3015:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(15));
	CUT_3016:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(16));
	CUT_3017:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(17));
	CUT_3018:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(18));
	CUT_3019:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(19));
	CUT_3020:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(20));
	CUT_3021:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(21));
	CUT_3022:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(22));
	CUT_3023:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(23));
	CUT_3024:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(24));
	CUT_3025:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(25));
	CUT_3026:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(26));
	CUT_3027:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(27));
	CUT_3028:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(28));
	CUT_3029:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(29));
	CUT_3030:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(30));
	CUT_3031:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(31));
	CUT_3032:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(32));
	CUT_3033:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(33));
	CUT_3034:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(34));
	CUT_3035:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(35));
	CUT_3036:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(36));
	CUT_3037:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(37));
	CUT_3038:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(38));
	CUT_3039:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(39));
	CUT_3040:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(40));
	CUT_3041:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(41));
	CUT_3042:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(42));
	CUT_3043:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(43));
	CUT_3044:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(44));
	CUT_3045:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(45));
	CUT_3046:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(46));
	CUT_3047:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(47));
	CUT_3048:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(48));
	CUT_3049:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(60)(49));
	CUT_3050:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(0));
	CUT_3051:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(1));
	CUT_3052:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(2));
	CUT_3053:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(3));
	CUT_3054:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(4));
	CUT_3055:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(5));
	CUT_3056:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(6));
	CUT_3057:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(7));
	CUT_3058:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(8));
	CUT_3059:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(9));
	CUT_3060:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(10));
	CUT_3061:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(11));
	CUT_3062:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(12));
	CUT_3063:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(13));
	CUT_3064:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(14));
	CUT_3065:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(15));
	CUT_3066:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(16));
	CUT_3067:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(17));
	CUT_3068:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(18));
	CUT_3069:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(19));
	CUT_3070:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(20));
	CUT_3071:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(21));
	CUT_3072:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(22));
	CUT_3073:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(23));
	CUT_3074:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(24));
	CUT_3075:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(25));
	CUT_3076:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(26));
	CUT_3077:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(27));
	CUT_3078:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(28));
	CUT_3079:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(29));
	CUT_3080:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(30));
	CUT_3081:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(31));
	CUT_3082:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(32));
	CUT_3083:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(33));
	CUT_3084:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(34));
	CUT_3085:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(35));
	CUT_3086:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(36));
	CUT_3087:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(37));
	CUT_3088:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(38));
	CUT_3089:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(39));
	CUT_3090:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(40));
	CUT_3091:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(41));
	CUT_3092:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(42));
	CUT_3093:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(43));
	CUT_3094:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(44));
	CUT_3095:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(45));
	CUT_3096:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(46));
	CUT_3097:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(47));
	CUT_3098:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(48));
	CUT_3099:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(61)(49));
	CUT_3100:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(0));
	CUT_3101:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(1));
	CUT_3102:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(2));
	CUT_3103:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(3));
	CUT_3104:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(4));
	CUT_3105:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(5));
	CUT_3106:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(6));
	CUT_3107:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(7));
	CUT_3108:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(8));
	CUT_3109:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(9));
	CUT_3110:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(10));
	CUT_3111:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(11));
	CUT_3112:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(12));
	CUT_3113:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(13));
	CUT_3114:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(14));
	CUT_3115:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(15));
	CUT_3116:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(16));
	CUT_3117:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(17));
	CUT_3118:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(18));
	CUT_3119:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(19));
	CUT_3120:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(20));
	CUT_3121:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(21));
	CUT_3122:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(22));
	CUT_3123:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(23));
	CUT_3124:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(24));
	CUT_3125:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(25));
	CUT_3126:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(26));
	CUT_3127:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(27));
	CUT_3128:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(28));
	CUT_3129:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(29));
	CUT_3130:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(30));
	CUT_3131:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(31));
	CUT_3132:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(32));
	CUT_3133:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(33));
	CUT_3134:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(34));
	CUT_3135:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(35));
	CUT_3136:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(36));
	CUT_3137:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(37));
	CUT_3138:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(38));
	CUT_3139:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(39));
	CUT_3140:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(40));
	CUT_3141:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(41));
	CUT_3142:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(42));
	CUT_3143:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(43));
	CUT_3144:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(44));
	CUT_3145:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(45));
	CUT_3146:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(46));
	CUT_3147:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(47));
	CUT_3148:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(48));
	CUT_3149:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(62)(49));
	CUT_3150:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(0));
	CUT_3151:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(1));
	CUT_3152:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(2));
	CUT_3153:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(3));
	CUT_3154:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(4));
	CUT_3155:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(5));
	CUT_3156:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(6));
	CUT_3157:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(7));
	CUT_3158:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(8));
	CUT_3159:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(9));
	CUT_3160:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(10));
	CUT_3161:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(11));
	CUT_3162:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(12));
	CUT_3163:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(13));
	CUT_3164:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(14));
	CUT_3165:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(15));
	CUT_3166:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(16));
	CUT_3167:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(17));
	CUT_3168:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(18));
	CUT_3169:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(19));
	CUT_3170:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(20));
	CUT_3171:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(21));
	CUT_3172:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(22));
	CUT_3173:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(23));
	CUT_3174:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(24));
	CUT_3175:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(25));
	CUT_3176:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(26));
	CUT_3177:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(27));
	CUT_3178:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(28));
	CUT_3179:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(29));
	CUT_3180:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(30));
	CUT_3181:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(31));
	CUT_3182:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(32));
	CUT_3183:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(33));
	CUT_3184:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(34));
	CUT_3185:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(35));
	CUT_3186:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(36));
	CUT_3187:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(37));
	CUT_3188:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(38));
	CUT_3189:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(39));
	CUT_3190:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(40));
	CUT_3191:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(41));
	CUT_3192:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(42));
	CUT_3193:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(43));
	CUT_3194:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(44));
	CUT_3195:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(45));
	CUT_3196:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(46));
	CUT_3197:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(47));
	CUT_3198:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(48));
	CUT_3199:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(63)(49));
	CUT_3200:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(0));
	CUT_3201:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(1));
	CUT_3202:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(2));
	CUT_3203:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(3));
	CUT_3204:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(4));
	CUT_3205:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(5));
	CUT_3206:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(6));
	CUT_3207:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(7));
	CUT_3208:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(8));
	CUT_3209:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(9));
	CUT_3210:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(10));
	CUT_3211:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(11));
	CUT_3212:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(12));
	CUT_3213:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(13));
	CUT_3214:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(14));
	CUT_3215:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(15));
	CUT_3216:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(16));
	CUT_3217:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(17));
	CUT_3218:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(18));
	CUT_3219:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(19));
	CUT_3220:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(20));
	CUT_3221:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(21));
	CUT_3222:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(22));
	CUT_3223:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(23));
	CUT_3224:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(24));
	CUT_3225:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(25));
	CUT_3226:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(26));
	CUT_3227:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(27));
	CUT_3228:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(28));
	CUT_3229:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(29));
	CUT_3230:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(30));
	CUT_3231:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(31));
	CUT_3232:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(32));
	CUT_3233:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(33));
	CUT_3234:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(34));
	CUT_3235:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(35));
	CUT_3236:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(36));
	CUT_3237:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(37));
	CUT_3238:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(38));
	CUT_3239:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(39));
	CUT_3240:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(40));
	CUT_3241:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(41));
	CUT_3242:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(42));
	CUT_3243:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(43));
	CUT_3244:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(44));
	CUT_3245:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(45));
	CUT_3246:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(46));
	CUT_3247:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(47));
	CUT_3248:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(48));
	CUT_3249:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(64)(49));
	CUT_3250:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(0));
	CUT_3251:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(1));
	CUT_3252:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(2));
	CUT_3253:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(3));
	CUT_3254:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(4));
	CUT_3255:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(5));
	CUT_3256:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(6));
	CUT_3257:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(7));
	CUT_3258:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(8));
	CUT_3259:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(9));
	CUT_3260:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(10));
	CUT_3261:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(11));
	CUT_3262:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(12));
	CUT_3263:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(13));
	CUT_3264:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(14));
	CUT_3265:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(15));
	CUT_3266:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(16));
	CUT_3267:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(17));
	CUT_3268:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(18));
	CUT_3269:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(19));
	CUT_3270:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(20));
	CUT_3271:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(21));
	CUT_3272:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(22));
	CUT_3273:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(23));
	CUT_3274:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(24));
	CUT_3275:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(25));
	CUT_3276:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(26));
	CUT_3277:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(27));
	CUT_3278:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(28));
	CUT_3279:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(29));
	CUT_3280:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(30));
	CUT_3281:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(31));
	CUT_3282:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(32));
	CUT_3283:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(33));
	CUT_3284:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(34));
	CUT_3285:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(35));
	CUT_3286:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(36));
	CUT_3287:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(37));
	CUT_3288:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(38));
	CUT_3289:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(39));
	CUT_3290:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(40));
	CUT_3291:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(41));
	CUT_3292:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(42));
	CUT_3293:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(43));
	CUT_3294:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(44));
	CUT_3295:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(45));
	CUT_3296:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(46));
	CUT_3297:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(47));
	CUT_3298:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(48));
	CUT_3299:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(65)(49));
	CUT_3300:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(0));
	CUT_3301:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(1));
	CUT_3302:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(2));
	CUT_3303:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(3));
	CUT_3304:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(4));
	CUT_3305:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(5));
	CUT_3306:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(6));
	CUT_3307:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(7));
	CUT_3308:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(8));
	CUT_3309:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(9));
	CUT_3310:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(10));
	CUT_3311:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(11));
	CUT_3312:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(12));
	CUT_3313:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(13));
	CUT_3314:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(14));
	CUT_3315:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(15));
	CUT_3316:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(16));
	CUT_3317:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(17));
	CUT_3318:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(18));
	CUT_3319:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(19));
	CUT_3320:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(20));
	CUT_3321:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(21));
	CUT_3322:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(22));
	CUT_3323:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(23));
	CUT_3324:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(24));
	CUT_3325:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(25));
	CUT_3326:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(26));
	CUT_3327:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(27));
	CUT_3328:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(28));
	CUT_3329:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(29));
	CUT_3330:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(30));
	CUT_3331:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(31));
	CUT_3332:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(32));
	CUT_3333:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(33));
	CUT_3334:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(34));
	CUT_3335:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(35));
	CUT_3336:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(36));
	CUT_3337:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(37));
	CUT_3338:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(38));
	CUT_3339:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(39));
	CUT_3340:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(40));
	CUT_3341:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(41));
	CUT_3342:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(42));
	CUT_3343:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(43));
	CUT_3344:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(44));
	CUT_3345:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(45));
	CUT_3346:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(46));
	CUT_3347:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(47));
	CUT_3348:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(48));
	CUT_3349:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(66)(49));
	CUT_3350:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(0));
	CUT_3351:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(1));
	CUT_3352:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(2));
	CUT_3353:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(3));
	CUT_3354:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(4));
	CUT_3355:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(5));
	CUT_3356:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(6));
	CUT_3357:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(7));
	CUT_3358:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(8));
	CUT_3359:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(9));
	CUT_3360:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(10));
	CUT_3361:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(11));
	CUT_3362:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(12));
	CUT_3363:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(13));
	CUT_3364:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(14));
	CUT_3365:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(15));
	CUT_3366:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(16));
	CUT_3367:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(17));
	CUT_3368:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(18));
	CUT_3369:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(19));
	CUT_3370:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(20));
	CUT_3371:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(21));
	CUT_3372:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(22));
	CUT_3373:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(23));
	CUT_3374:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(24));
	CUT_3375:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(25));
	CUT_3376:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(26));
	CUT_3377:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(27));
	CUT_3378:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(28));
	CUT_3379:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(29));
	CUT_3380:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(30));
	CUT_3381:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(31));
	CUT_3382:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(32));
	CUT_3383:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(33));
	CUT_3384:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(34));
	CUT_3385:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(35));
	CUT_3386:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(36));
	CUT_3387:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(37));
	CUT_3388:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(38));
	CUT_3389:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(39));
	CUT_3390:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(40));
	CUT_3391:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(41));
	CUT_3392:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(42));
	CUT_3393:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(43));
	CUT_3394:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(44));
	CUT_3395:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(45));
	CUT_3396:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(46));
	CUT_3397:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(47));
	CUT_3398:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(48));
	CUT_3399:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(67)(49));
	CUT_3400:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(0));
	CUT_3401:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(1));
	CUT_3402:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(2));
	CUT_3403:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(3));
	CUT_3404:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(4));
	CUT_3405:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(5));
	CUT_3406:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(6));
	CUT_3407:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(7));
	CUT_3408:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(8));
	CUT_3409:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(9));
	CUT_3410:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(10));
	CUT_3411:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(11));
	CUT_3412:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(12));
	CUT_3413:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(13));
	CUT_3414:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(14));
	CUT_3415:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(15));
	CUT_3416:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(16));
	CUT_3417:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(17));
	CUT_3418:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(18));
	CUT_3419:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(19));
	CUT_3420:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(20));
	CUT_3421:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(21));
	CUT_3422:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(22));
	CUT_3423:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(23));
	CUT_3424:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(24));
	CUT_3425:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(25));
	CUT_3426:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(26));
	CUT_3427:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(27));
	CUT_3428:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(28));
	CUT_3429:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(29));
	CUT_3430:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(30));
	CUT_3431:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(31));
	CUT_3432:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(32));
	CUT_3433:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(33));
	CUT_3434:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(34));
	CUT_3435:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(35));
	CUT_3436:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(36));
	CUT_3437:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(37));
	CUT_3438:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(38));
	CUT_3439:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(39));
	CUT_3440:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(40));
	CUT_3441:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(41));
	CUT_3442:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(42));
	CUT_3443:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(43));
	CUT_3444:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(44));
	CUT_3445:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(45));
	CUT_3446:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(46));
	CUT_3447:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(47));
	CUT_3448:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(48));
	CUT_3449:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(68)(49));
	CUT_3450:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(0));
	CUT_3451:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(1));
	CUT_3452:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(2));
	CUT_3453:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(3));
	CUT_3454:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(4));
	CUT_3455:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(5));
	CUT_3456:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(6));
	CUT_3457:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(7));
	CUT_3458:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(8));
	CUT_3459:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(9));
	CUT_3460:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(10));
	CUT_3461:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(11));
	CUT_3462:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(12));
	CUT_3463:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(13));
	CUT_3464:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(14));
	CUT_3465:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(15));
	CUT_3466:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(16));
	CUT_3467:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(17));
	CUT_3468:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(18));
	CUT_3469:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(19));
	CUT_3470:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(20));
	CUT_3471:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(21));
	CUT_3472:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(22));
	CUT_3473:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(23));
	CUT_3474:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(24));
	CUT_3475:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(25));
	CUT_3476:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(26));
	CUT_3477:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(27));
	CUT_3478:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(28));
	CUT_3479:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(29));
	CUT_3480:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(30));
	CUT_3481:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(31));
	CUT_3482:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(32));
	CUT_3483:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(33));
	CUT_3484:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(34));
	CUT_3485:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(35));
	CUT_3486:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(36));
	CUT_3487:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(37));
	CUT_3488:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(38));
	CUT_3489:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(39));
	CUT_3490:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(40));
	CUT_3491:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(41));
	CUT_3492:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(42));
	CUT_3493:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(43));
	CUT_3494:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(44));
	CUT_3495:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(45));
	CUT_3496:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(46));
	CUT_3497:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(47));
	CUT_3498:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(48));
	CUT_3499:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(69)(49));
	CUT_3500:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(0));
	CUT_3501:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(1));
	CUT_3502:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(2));
	CUT_3503:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(3));
	CUT_3504:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(4));
	CUT_3505:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(5));
	CUT_3506:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(6));
	CUT_3507:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(7));
	CUT_3508:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(8));
	CUT_3509:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(9));
	CUT_3510:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(10));
	CUT_3511:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(11));
	CUT_3512:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(12));
	CUT_3513:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(13));
	CUT_3514:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(14));
	CUT_3515:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(15));
	CUT_3516:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(16));
	CUT_3517:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(17));
	CUT_3518:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(18));
	CUT_3519:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(19));
	CUT_3520:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(20));
	CUT_3521:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(21));
	CUT_3522:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(22));
	CUT_3523:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(23));
	CUT_3524:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(24));
	CUT_3525:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(25));
	CUT_3526:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(26));
	CUT_3527:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(27));
	CUT_3528:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(28));
	CUT_3529:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(29));
	CUT_3530:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(30));
	CUT_3531:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(31));
	CUT_3532:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(32));
	CUT_3533:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(33));
	CUT_3534:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(34));
	CUT_3535:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(35));
	CUT_3536:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(36));
	CUT_3537:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(37));
	CUT_3538:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(38));
	CUT_3539:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(39));
	CUT_3540:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(40));
	CUT_3541:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(41));
	CUT_3542:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(42));
	CUT_3543:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(43));
	CUT_3544:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(44));
	CUT_3545:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(45));
	CUT_3546:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(46));
	CUT_3547:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(47));
	CUT_3548:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(48));
	CUT_3549:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(70)(49));
	CUT_3550:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(0));
	CUT_3551:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(1));
	CUT_3552:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(2));
	CUT_3553:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(3));
	CUT_3554:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(4));
	CUT_3555:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(5));
	CUT_3556:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(6));
	CUT_3557:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(7));
	CUT_3558:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(8));
	CUT_3559:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(9));
	CUT_3560:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(10));
	CUT_3561:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(11));
	CUT_3562:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(12));
	CUT_3563:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(13));
	CUT_3564:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(14));
	CUT_3565:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(15));
	CUT_3566:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(16));
	CUT_3567:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(17));
	CUT_3568:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(18));
	CUT_3569:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(19));
	CUT_3570:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(20));
	CUT_3571:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(21));
	CUT_3572:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(22));
	CUT_3573:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(23));
	CUT_3574:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(24));
	CUT_3575:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(25));
	CUT_3576:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(26));
	CUT_3577:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(27));
	CUT_3578:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(28));
	CUT_3579:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(29));
	CUT_3580:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(30));
	CUT_3581:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(31));
	CUT_3582:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(32));
	CUT_3583:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(33));
	CUT_3584:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(34));
	CUT_3585:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(35));
	CUT_3586:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(36));
	CUT_3587:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(37));
	CUT_3588:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(38));
	CUT_3589:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(39));
	CUT_3590:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(40));
	CUT_3591:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(41));
	CUT_3592:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(42));
	CUT_3593:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(43));
	CUT_3594:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(44));
	CUT_3595:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(45));
	CUT_3596:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(46));
	CUT_3597:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(47));
	CUT_3598:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(48));
	CUT_3599:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(71)(49));
	CUT_3600:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(0));
	CUT_3601:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(1));
	CUT_3602:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(2));
	CUT_3603:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(3));
	CUT_3604:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(4));
	CUT_3605:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(5));
	CUT_3606:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(6));
	CUT_3607:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(7));
	CUT_3608:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(8));
	CUT_3609:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(9));
	CUT_3610:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(10));
	CUT_3611:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(11));
	CUT_3612:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(12));
	CUT_3613:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(13));
	CUT_3614:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(14));
	CUT_3615:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(15));
	CUT_3616:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(16));
	CUT_3617:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(17));
	CUT_3618:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(18));
	CUT_3619:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(19));
	CUT_3620:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(20));
	CUT_3621:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(21));
	CUT_3622:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(22));
	CUT_3623:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(23));
	CUT_3624:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(24));
	CUT_3625:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(25));
	CUT_3626:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(26));
	CUT_3627:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(27));
	CUT_3628:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(28));
	CUT_3629:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(29));
	CUT_3630:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(30));
	CUT_3631:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(31));
	CUT_3632:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(32));
	CUT_3633:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(33));
	CUT_3634:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(34));
	CUT_3635:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(35));
	CUT_3636:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(36));
	CUT_3637:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(37));
	CUT_3638:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(38));
	CUT_3639:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(39));
	CUT_3640:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(40));
	CUT_3641:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(41));
	CUT_3642:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(42));
	CUT_3643:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(43));
	CUT_3644:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(44));
	CUT_3645:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(45));
	CUT_3646:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(46));
	CUT_3647:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(47));
	CUT_3648:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(48));
	CUT_3649:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(72)(49));
	CUT_3650:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(0));
	CUT_3651:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(1));
	CUT_3652:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(2));
	CUT_3653:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(3));
	CUT_3654:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(4));
	CUT_3655:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(5));
	CUT_3656:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(6));
	CUT_3657:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(7));
	CUT_3658:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(8));
	CUT_3659:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(9));
	CUT_3660:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(10));
	CUT_3661:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(11));
	CUT_3662:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(12));
	CUT_3663:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(13));
	CUT_3664:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(14));
	CUT_3665:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(15));
	CUT_3666:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(16));
	CUT_3667:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(17));
	CUT_3668:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(18));
	CUT_3669:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(19));
	CUT_3670:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(20));
	CUT_3671:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(21));
	CUT_3672:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(22));
	CUT_3673:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(23));
	CUT_3674:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(24));
	CUT_3675:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(25));
	CUT_3676:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(26));
	CUT_3677:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(27));
	CUT_3678:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(28));
	CUT_3679:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(29));
	CUT_3680:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(30));
	CUT_3681:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(31));
	CUT_3682:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(32));
	CUT_3683:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(33));
	CUT_3684:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(34));
	CUT_3685:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(35));
	CUT_3686:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(36));
	CUT_3687:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(37));
	CUT_3688:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(38));
	CUT_3689:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(39));
	CUT_3690:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(40));
	CUT_3691:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(41));
	CUT_3692:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(42));
	CUT_3693:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(43));
	CUT_3694:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(44));
	CUT_3695:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(45));
	CUT_3696:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(46));
	CUT_3697:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(47));
	CUT_3698:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(48));
	CUT_3699:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(73)(49));
	CUT_3700:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(0));
	CUT_3701:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(1));
	CUT_3702:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(2));
	CUT_3703:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(3));
	CUT_3704:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(4));
	CUT_3705:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(5));
	CUT_3706:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(6));
	CUT_3707:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(7));
	CUT_3708:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(8));
	CUT_3709:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(9));
	CUT_3710:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(10));
	CUT_3711:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(11));
	CUT_3712:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(12));
	CUT_3713:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(13));
	CUT_3714:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(14));
	CUT_3715:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(15));
	CUT_3716:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(16));
	CUT_3717:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(17));
	CUT_3718:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(18));
	CUT_3719:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(19));
	CUT_3720:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(20));
	CUT_3721:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(21));
	CUT_3722:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(22));
	CUT_3723:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(23));
	CUT_3724:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(24));
	CUT_3725:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(25));
	CUT_3726:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(26));
	CUT_3727:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(27));
	CUT_3728:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(28));
	CUT_3729:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(29));
	CUT_3730:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(30));
	CUT_3731:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(31));
	CUT_3732:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(32));
	CUT_3733:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(33));
	CUT_3734:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(34));
	CUT_3735:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(35));
	CUT_3736:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(36));
	CUT_3737:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(37));
	CUT_3738:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(38));
	CUT_3739:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(39));
	CUT_3740:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(40));
	CUT_3741:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(41));
	CUT_3742:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(42));
	CUT_3743:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(43));
	CUT_3744:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(44));
	CUT_3745:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(45));
	CUT_3746:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(46));
	CUT_3747:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(47));
	CUT_3748:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(48));
	CUT_3749:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(74)(49));
	CUT_3750:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(0));
	CUT_3751:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(1));
	CUT_3752:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(2));
	CUT_3753:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(3));
	CUT_3754:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(4));
	CUT_3755:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(5));
	CUT_3756:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(6));
	CUT_3757:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(7));
	CUT_3758:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(8));
	CUT_3759:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(9));
	CUT_3760:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(10));
	CUT_3761:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(11));
	CUT_3762:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(12));
	CUT_3763:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(13));
	CUT_3764:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(14));
	CUT_3765:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(15));
	CUT_3766:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(16));
	CUT_3767:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(17));
	CUT_3768:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(18));
	CUT_3769:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(19));
	CUT_3770:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(20));
	CUT_3771:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(21));
	CUT_3772:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(22));
	CUT_3773:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(23));
	CUT_3774:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(24));
	CUT_3775:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(25));
	CUT_3776:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(26));
	CUT_3777:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(27));
	CUT_3778:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(28));
	CUT_3779:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(29));
	CUT_3780:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(30));
	CUT_3781:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(31));
	CUT_3782:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(32));
	CUT_3783:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(33));
	CUT_3784:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(34));
	CUT_3785:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(35));
	CUT_3786:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(36));
	CUT_3787:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(37));
	CUT_3788:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(38));
	CUT_3789:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(39));
	CUT_3790:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(40));
	CUT_3791:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(41));
	CUT_3792:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(42));
	CUT_3793:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(43));
	CUT_3794:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(44));
	CUT_3795:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(45));
	CUT_3796:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(46));
	CUT_3797:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(47));
	CUT_3798:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(48));
	CUT_3799:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(75)(49));
	CUT_3800:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(0));
	CUT_3801:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(1));
	CUT_3802:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(2));
	CUT_3803:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(3));
	CUT_3804:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(4));
	CUT_3805:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(5));
	CUT_3806:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(6));
	CUT_3807:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(7));
	CUT_3808:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(8));
	CUT_3809:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(9));
	CUT_3810:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(10));
	CUT_3811:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(11));
	CUT_3812:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(12));
	CUT_3813:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(13));
	CUT_3814:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(14));
	CUT_3815:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(15));
	CUT_3816:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(16));
	CUT_3817:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(17));
	CUT_3818:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(18));
	CUT_3819:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(19));
	CUT_3820:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(20));
	CUT_3821:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(21));
	CUT_3822:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(22));
	CUT_3823:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(23));
	CUT_3824:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(24));
	CUT_3825:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(25));
	CUT_3826:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(26));
	CUT_3827:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(27));
	CUT_3828:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(28));
	CUT_3829:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(29));
	CUT_3830:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(30));
	CUT_3831:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(31));
	CUT_3832:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(32));
	CUT_3833:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(33));
	CUT_3834:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(34));
	CUT_3835:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(35));
	CUT_3836:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(36));
	CUT_3837:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(37));
	CUT_3838:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(38));
	CUT_3839:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(39));
	CUT_3840:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(40));
	CUT_3841:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(41));
	CUT_3842:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(42));
	CUT_3843:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(43));
	CUT_3844:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(44));
	CUT_3845:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(45));
	CUT_3846:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(46));
	CUT_3847:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(47));
	CUT_3848:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(48));
	CUT_3849:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(76)(49));
	CUT_3850:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(0));
	CUT_3851:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(1));
	CUT_3852:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(2));
	CUT_3853:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(3));
	CUT_3854:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(4));
	CUT_3855:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(5));
	CUT_3856:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(6));
	CUT_3857:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(7));
	CUT_3858:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(8));
	CUT_3859:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(9));
	CUT_3860:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(10));
	CUT_3861:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(11));
	CUT_3862:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(12));
	CUT_3863:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(13));
	CUT_3864:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(14));
	CUT_3865:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(15));
	CUT_3866:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(16));
	CUT_3867:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(17));
	CUT_3868:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(18));
	CUT_3869:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(19));
	CUT_3870:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(20));
	CUT_3871:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(21));
	CUT_3872:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(22));
	CUT_3873:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(23));
	CUT_3874:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(24));
	CUT_3875:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(25));
	CUT_3876:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(26));
	CUT_3877:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(27));
	CUT_3878:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(28));
	CUT_3879:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(29));
	CUT_3880:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(30));
	CUT_3881:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(31));
	CUT_3882:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(32));
	CUT_3883:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(33));
	CUT_3884:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(34));
	CUT_3885:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(35));
	CUT_3886:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(36));
	CUT_3887:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(37));
	CUT_3888:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(38));
	CUT_3889:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(39));
	CUT_3890:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(40));
	CUT_3891:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(41));
	CUT_3892:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(42));
	CUT_3893:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(43));
	CUT_3894:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(44));
	CUT_3895:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(45));
	CUT_3896:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(46));
	CUT_3897:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(47));
	CUT_3898:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(48));
	CUT_3899:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(77)(49));
	CUT_3900:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(0));
	CUT_3901:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(1));
	CUT_3902:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(2));
	CUT_3903:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(3));
	CUT_3904:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(4));
	CUT_3905:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(5));
	CUT_3906:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(6));
	CUT_3907:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(7));
	CUT_3908:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(8));
	CUT_3909:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(9));
	CUT_3910:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(10));
	CUT_3911:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(11));
	CUT_3912:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(12));
	CUT_3913:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(13));
	CUT_3914:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(14));
	CUT_3915:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(15));
	CUT_3916:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(16));
	CUT_3917:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(17));
	CUT_3918:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(18));
	CUT_3919:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(19));
	CUT_3920:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(20));
	CUT_3921:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(21));
	CUT_3922:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(22));
	CUT_3923:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(23));
	CUT_3924:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(24));
	CUT_3925:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(25));
	CUT_3926:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(26));
	CUT_3927:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(27));
	CUT_3928:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(28));
	CUT_3929:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(29));
	CUT_3930:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(30));
	CUT_3931:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(31));
	CUT_3932:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(32));
	CUT_3933:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(33));
	CUT_3934:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(34));
	CUT_3935:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(35));
	CUT_3936:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(36));
	CUT_3937:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(37));
	CUT_3938:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(38));
	CUT_3939:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(39));
	CUT_3940:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(40));
	CUT_3941:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(41));
	CUT_3942:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(42));
	CUT_3943:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(43));
	CUT_3944:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(44));
	CUT_3945:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(45));
	CUT_3946:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(46));
	CUT_3947:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(47));
	CUT_3948:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(48));
	CUT_3949:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(78)(49));
	CUT_3950:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(0));
	CUT_3951:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(1));
	CUT_3952:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(2));
	CUT_3953:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(3));
	CUT_3954:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(4));
	CUT_3955:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(5));
	CUT_3956:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(6));
	CUT_3957:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(7));
	CUT_3958:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(8));
	CUT_3959:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(9));
	CUT_3960:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(10));
	CUT_3961:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(11));
	CUT_3962:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(12));
	CUT_3963:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(13));
	CUT_3964:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(14));
	CUT_3965:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(15));
	CUT_3966:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(16));
	CUT_3967:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(17));
	CUT_3968:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(18));
	CUT_3969:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(19));
	CUT_3970:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(20));
	CUT_3971:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(21));
	CUT_3972:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(22));
	CUT_3973:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(23));
	CUT_3974:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(24));
	CUT_3975:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(25));
	CUT_3976:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(26));
	CUT_3977:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(27));
	CUT_3978:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(28));
	CUT_3979:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(29));
	CUT_3980:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(30));
	CUT_3981:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(31));
	CUT_3982:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(32));
	CUT_3983:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(33));
	CUT_3984:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(34));
	CUT_3985:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(35));
	CUT_3986:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(36));
	CUT_3987:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(37));
	CUT_3988:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(38));
	CUT_3989:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(39));
	CUT_3990:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(40));
	CUT_3991:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(41));
	CUT_3992:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(42));
	CUT_3993:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(43));
	CUT_3994:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(44));
	CUT_3995:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(45));
	CUT_3996:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(46));
	CUT_3997:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(47));
	CUT_3998:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(48));
	CUT_3999:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(79)(49));
	CUT_4000:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(0));
	CUT_4001:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(1));
	CUT_4002:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(2));
	CUT_4003:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(3));
	CUT_4004:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(4));
	CUT_4005:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(5));
	CUT_4006:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(6));
	CUT_4007:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(7));
	CUT_4008:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(8));
	CUT_4009:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(9));
	CUT_4010:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(10));
	CUT_4011:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(11));
	CUT_4012:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(12));
	CUT_4013:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(13));
	CUT_4014:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(14));
	CUT_4015:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(15));
	CUT_4016:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(16));
	CUT_4017:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(17));
	CUT_4018:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(18));
	CUT_4019:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(19));
	CUT_4020:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(20));
	CUT_4021:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(21));
	CUT_4022:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(22));
	CUT_4023:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(23));
	CUT_4024:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(24));
	CUT_4025:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(25));
	CUT_4026:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(26));
	CUT_4027:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(27));
	CUT_4028:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(28));
	CUT_4029:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(29));
	CUT_4030:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(30));
	CUT_4031:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(31));
	CUT_4032:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(32));
	CUT_4033:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(33));
	CUT_4034:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(34));
	CUT_4035:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(35));
	CUT_4036:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(36));
	CUT_4037:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(37));
	CUT_4038:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(38));
	CUT_4039:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(39));
	CUT_4040:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(40));
	CUT_4041:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(41));
	CUT_4042:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(42));
	CUT_4043:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(43));
	CUT_4044:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(44));
	CUT_4045:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(45));
	CUT_4046:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(46));
	CUT_4047:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(47));
	CUT_4048:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(48));
	CUT_4049:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(80)(49));
	CUT_4050:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(0));
	CUT_4051:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(1));
	CUT_4052:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(2));
	CUT_4053:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(3));
	CUT_4054:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(4));
	CUT_4055:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(5));
	CUT_4056:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(6));
	CUT_4057:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(7));
	CUT_4058:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(8));
	CUT_4059:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(9));
	CUT_4060:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(10));
	CUT_4061:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(11));
	CUT_4062:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(12));
	CUT_4063:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(13));
	CUT_4064:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(14));
	CUT_4065:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(15));
	CUT_4066:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(16));
	CUT_4067:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(17));
	CUT_4068:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(18));
	CUT_4069:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(19));
	CUT_4070:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(20));
	CUT_4071:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(21));
	CUT_4072:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(22));
	CUT_4073:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(23));
	CUT_4074:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(24));
	CUT_4075:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(25));
	CUT_4076:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(26));
	CUT_4077:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(27));
	CUT_4078:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(28));
	CUT_4079:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(29));
	CUT_4080:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(30));
	CUT_4081:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(31));
	CUT_4082:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(32));
	CUT_4083:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(33));
	CUT_4084:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(34));
	CUT_4085:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(35));
	CUT_4086:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(36));
	CUT_4087:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(37));
	CUT_4088:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(38));
	CUT_4089:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(39));
	CUT_4090:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(40));
	CUT_4091:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(41));
	CUT_4092:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(42));
	CUT_4093:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(43));
	CUT_4094:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(44));
	CUT_4095:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(45));
	CUT_4096:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(46));
	CUT_4097:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(47));
	CUT_4098:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(48));
	CUT_4099:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(81)(49));
	CUT_4100:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(0));
	CUT_4101:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(1));
	CUT_4102:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(2));
	CUT_4103:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(3));
	CUT_4104:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(4));
	CUT_4105:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(5));
	CUT_4106:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(6));
	CUT_4107:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(7));
	CUT_4108:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(8));
	CUT_4109:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(9));
	CUT_4110:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(10));
	CUT_4111:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(11));
	CUT_4112:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(12));
	CUT_4113:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(13));
	CUT_4114:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(14));
	CUT_4115:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(15));
	CUT_4116:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(16));
	CUT_4117:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(17));
	CUT_4118:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(18));
	CUT_4119:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(19));
	CUT_4120:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(20));
	CUT_4121:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(21));
	CUT_4122:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(22));
	CUT_4123:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(23));
	CUT_4124:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(24));
	CUT_4125:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(25));
	CUT_4126:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(26));
	CUT_4127:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(27));
	CUT_4128:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(28));
	CUT_4129:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(29));
	CUT_4130:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(30));
	CUT_4131:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(31));
	CUT_4132:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(32));
	CUT_4133:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(33));
	CUT_4134:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(34));
	CUT_4135:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(35));
	CUT_4136:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(36));
	CUT_4137:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(37));
	CUT_4138:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(38));
	CUT_4139:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(39));
	CUT_4140:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(40));
	CUT_4141:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(41));
	CUT_4142:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(42));
	CUT_4143:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(43));
	CUT_4144:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(44));
	CUT_4145:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(45));
	CUT_4146:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(46));
	CUT_4147:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(47));
	CUT_4148:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(48));
	CUT_4149:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(82)(49));
	CUT_4150:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(0));
	CUT_4151:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(1));
	CUT_4152:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(2));
	CUT_4153:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(3));
	CUT_4154:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(4));
	CUT_4155:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(5));
	CUT_4156:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(6));
	CUT_4157:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(7));
	CUT_4158:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(8));
	CUT_4159:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(9));
	CUT_4160:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(10));
	CUT_4161:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(11));
	CUT_4162:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(12));
	CUT_4163:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(13));
	CUT_4164:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(14));
	CUT_4165:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(15));
	CUT_4166:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(16));
	CUT_4167:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(17));
	CUT_4168:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(18));
	CUT_4169:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(19));
	CUT_4170:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(20));
	CUT_4171:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(21));
	CUT_4172:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(22));
	CUT_4173:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(23));
	CUT_4174:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(24));
	CUT_4175:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(25));
	CUT_4176:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(26));
	CUT_4177:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(27));
	CUT_4178:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(28));
	CUT_4179:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(29));
	CUT_4180:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(30));
	CUT_4181:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(31));
	CUT_4182:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(32));
	CUT_4183:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(33));
	CUT_4184:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(34));
	CUT_4185:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(35));
	CUT_4186:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(36));
	CUT_4187:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(37));
	CUT_4188:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(38));
	CUT_4189:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(39));
	CUT_4190:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(40));
	CUT_4191:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(41));
	CUT_4192:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(42));
	CUT_4193:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(43));
	CUT_4194:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(44));
	CUT_4195:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(45));
	CUT_4196:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(46));
	CUT_4197:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(47));
	CUT_4198:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(48));
	CUT_4199:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(83)(49));
	CUT_4200:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(0));
	CUT_4201:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(1));
	CUT_4202:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(2));
	CUT_4203:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(3));
	CUT_4204:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(4));
	CUT_4205:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(5));
	CUT_4206:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(6));
	CUT_4207:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(7));
	CUT_4208:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(8));
	CUT_4209:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(9));
	CUT_4210:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(10));
	CUT_4211:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(11));
	CUT_4212:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(12));
	CUT_4213:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(13));
	CUT_4214:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(14));
	CUT_4215:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(15));
	CUT_4216:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(16));
	CUT_4217:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(17));
	CUT_4218:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(18));
	CUT_4219:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(19));
	CUT_4220:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(20));
	CUT_4221:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(21));
	CUT_4222:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(22));
	CUT_4223:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(23));
	CUT_4224:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(24));
	CUT_4225:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(25));
	CUT_4226:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(26));
	CUT_4227:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(27));
	CUT_4228:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(28));
	CUT_4229:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(29));
	CUT_4230:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(30));
	CUT_4231:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(31));
	CUT_4232:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(32));
	CUT_4233:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(33));
	CUT_4234:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(34));
	CUT_4235:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(35));
	CUT_4236:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(36));
	CUT_4237:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(37));
	CUT_4238:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(38));
	CUT_4239:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(39));
	CUT_4240:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(40));
	CUT_4241:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(41));
	CUT_4242:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(42));
	CUT_4243:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(43));
	CUT_4244:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(44));
	CUT_4245:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(45));
	CUT_4246:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(46));
	CUT_4247:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(47));
	CUT_4248:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(48));
	CUT_4249:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(84)(49));
	CUT_4250:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(0));
	CUT_4251:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(1));
	CUT_4252:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(2));
	CUT_4253:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(3));
	CUT_4254:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(4));
	CUT_4255:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(5));
	CUT_4256:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(6));
	CUT_4257:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(7));
	CUT_4258:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(8));
	CUT_4259:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(9));
	CUT_4260:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(10));
	CUT_4261:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(11));
	CUT_4262:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(12));
	CUT_4263:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(13));
	CUT_4264:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(14));
	CUT_4265:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(15));
	CUT_4266:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(16));
	CUT_4267:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(17));
	CUT_4268:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(18));
	CUT_4269:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(19));
	CUT_4270:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(20));
	CUT_4271:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(21));
	CUT_4272:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(22));
	CUT_4273:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(23));
	CUT_4274:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(24));
	CUT_4275:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(25));
	CUT_4276:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(26));
	CUT_4277:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(27));
	CUT_4278:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(28));
	CUT_4279:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(29));
	CUT_4280:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(30));
	CUT_4281:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(31));
	CUT_4282:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(32));
	CUT_4283:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(33));
	CUT_4284:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(34));
	CUT_4285:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(35));
	CUT_4286:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(36));
	CUT_4287:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(37));
	CUT_4288:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(38));
	CUT_4289:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(39));
	CUT_4290:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(40));
	CUT_4291:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(41));
	CUT_4292:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(42));
	CUT_4293:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(43));
	CUT_4294:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(44));
	CUT_4295:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(45));
	CUT_4296:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(46));
	CUT_4297:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(47));
	CUT_4298:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(48));
	CUT_4299:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(85)(49));
	CUT_4300:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(0));
	CUT_4301:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(1));
	CUT_4302:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(2));
	CUT_4303:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(3));
	CUT_4304:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(4));
	CUT_4305:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(5));
	CUT_4306:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(6));
	CUT_4307:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(7));
	CUT_4308:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(8));
	CUT_4309:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(9));
	CUT_4310:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(10));
	CUT_4311:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(11));
	CUT_4312:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(12));
	CUT_4313:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(13));
	CUT_4314:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(14));
	CUT_4315:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(15));
	CUT_4316:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(16));
	CUT_4317:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(17));
	CUT_4318:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(18));
	CUT_4319:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(19));
	CUT_4320:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(20));
	CUT_4321:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(21));
	CUT_4322:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(22));
	CUT_4323:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(23));
	CUT_4324:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(24));
	CUT_4325:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(25));
	CUT_4326:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(26));
	CUT_4327:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(27));
	CUT_4328:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(28));
	CUT_4329:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(29));
	CUT_4330:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(30));
	CUT_4331:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(31));
	CUT_4332:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(32));
	CUT_4333:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(33));
	CUT_4334:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(34));
	CUT_4335:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(35));
	CUT_4336:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(36));
	CUT_4337:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(37));
	CUT_4338:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(38));
	CUT_4339:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(39));
	CUT_4340:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(40));
	CUT_4341:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(41));
	CUT_4342:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(42));
	CUT_4343:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(43));
	CUT_4344:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(44));
	CUT_4345:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(45));
	CUT_4346:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(46));
	CUT_4347:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(47));
	CUT_4348:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(48));
	CUT_4349:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(86)(49));
	CUT_4350:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(0));
	CUT_4351:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(1));
	CUT_4352:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(2));
	CUT_4353:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(3));
	CUT_4354:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(4));
	CUT_4355:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(5));
	CUT_4356:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(6));
	CUT_4357:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(7));
	CUT_4358:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(8));
	CUT_4359:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(9));
	CUT_4360:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(10));
	CUT_4361:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(11));
	CUT_4362:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(12));
	CUT_4363:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(13));
	CUT_4364:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(14));
	CUT_4365:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(15));
	CUT_4366:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(16));
	CUT_4367:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(17));
	CUT_4368:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(18));
	CUT_4369:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(19));
	CUT_4370:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(20));
	CUT_4371:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(21));
	CUT_4372:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(22));
	CUT_4373:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(23));
	CUT_4374:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(24));
	CUT_4375:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(25));
	CUT_4376:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(26));
	CUT_4377:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(27));
	CUT_4378:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(28));
	CUT_4379:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(29));
	CUT_4380:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(30));
	CUT_4381:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(31));
	CUT_4382:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(32));
	CUT_4383:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(33));
	CUT_4384:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(34));
	CUT_4385:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(35));
	CUT_4386:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(36));
	CUT_4387:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(37));
	CUT_4388:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(38));
	CUT_4389:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(39));
	CUT_4390:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(40));
	CUT_4391:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(41));
	CUT_4392:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(42));
	CUT_4393:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(43));
	CUT_4394:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(44));
	CUT_4395:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(45));
	CUT_4396:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(46));
	CUT_4397:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(47));
	CUT_4398:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(48));
	CUT_4399:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(87)(49));
	CUT_4400:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(0));
	CUT_4401:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(1));
	CUT_4402:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(2));
	CUT_4403:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(3));
	CUT_4404:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(4));
	CUT_4405:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(5));
	CUT_4406:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(6));
	CUT_4407:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(7));
	CUT_4408:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(8));
	CUT_4409:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(9));
	CUT_4410:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(10));
	CUT_4411:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(11));
	CUT_4412:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(12));
	CUT_4413:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(13));
	CUT_4414:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(14));
	CUT_4415:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(15));
	CUT_4416:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(16));
	CUT_4417:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(17));
	CUT_4418:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(18));
	CUT_4419:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(19));
	CUT_4420:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(20));
	CUT_4421:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(21));
	CUT_4422:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(22));
	CUT_4423:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(23));
	CUT_4424:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(24));
	CUT_4425:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(25));
	CUT_4426:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(26));
	CUT_4427:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(27));
	CUT_4428:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(28));
	CUT_4429:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(29));
	CUT_4430:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(30));
	CUT_4431:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(31));
	CUT_4432:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(32));
	CUT_4433:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(33));
	CUT_4434:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(34));
	CUT_4435:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(35));
	CUT_4436:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(36));
	CUT_4437:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(37));
	CUT_4438:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(38));
	CUT_4439:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(39));
	CUT_4440:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(40));
	CUT_4441:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(41));
	CUT_4442:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(42));
	CUT_4443:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(43));
	CUT_4444:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(44));
	CUT_4445:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(45));
	CUT_4446:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(46));
	CUT_4447:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(47));
	CUT_4448:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(48));
	CUT_4449:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(88)(49));
	CUT_4450:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(0));
	CUT_4451:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(1));
	CUT_4452:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(2));
	CUT_4453:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(3));
	CUT_4454:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(4));
	CUT_4455:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(5));
	CUT_4456:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(6));
	CUT_4457:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(7));
	CUT_4458:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(8));
	CUT_4459:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(9));
	CUT_4460:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(10));
	CUT_4461:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(11));
	CUT_4462:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(12));
	CUT_4463:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(13));
	CUT_4464:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(14));
	CUT_4465:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(15));
	CUT_4466:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(16));
	CUT_4467:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(17));
	CUT_4468:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(18));
	CUT_4469:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(19));
	CUT_4470:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(20));
	CUT_4471:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(21));
	CUT_4472:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(22));
	CUT_4473:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(23));
	CUT_4474:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(24));
	CUT_4475:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(25));
	CUT_4476:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(26));
	CUT_4477:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(27));
	CUT_4478:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(28));
	CUT_4479:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(29));
	CUT_4480:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(30));
	CUT_4481:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(31));
	CUT_4482:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(32));
	CUT_4483:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(33));
	CUT_4484:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(34));
	CUT_4485:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(35));
	CUT_4486:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(36));
	CUT_4487:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(37));
	CUT_4488:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(38));
	CUT_4489:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(39));
	CUT_4490:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(40));
	CUT_4491:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(41));
	CUT_4492:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(42));
	CUT_4493:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(43));
	CUT_4494:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(44));
	CUT_4495:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(45));
	CUT_4496:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(46));
	CUT_4497:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(47));
	CUT_4498:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(48));
	CUT_4499:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(89)(49));
	CUT_4500:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(0));
	CUT_4501:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(1));
	CUT_4502:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(2));
	CUT_4503:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(3));
	CUT_4504:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(4));
	CUT_4505:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(5));
	CUT_4506:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(6));
	CUT_4507:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(7));
	CUT_4508:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(8));
	CUT_4509:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(9));
	CUT_4510:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(10));
	CUT_4511:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(11));
	CUT_4512:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(12));
	CUT_4513:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(13));
	CUT_4514:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(14));
	CUT_4515:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(15));
	CUT_4516:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(16));
	CUT_4517:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(17));
	CUT_4518:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(18));
	CUT_4519:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(19));
	CUT_4520:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(20));
	CUT_4521:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(21));
	CUT_4522:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(22));
	CUT_4523:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(23));
	CUT_4524:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(24));
	CUT_4525:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(25));
	CUT_4526:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(26));
	CUT_4527:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(27));
	CUT_4528:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(28));
	CUT_4529:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(29));
	CUT_4530:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(30));
	CUT_4531:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(31));
	CUT_4532:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(32));
	CUT_4533:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(33));
	CUT_4534:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(34));
	CUT_4535:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(35));
	CUT_4536:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(36));
	CUT_4537:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(37));
	CUT_4538:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(38));
	CUT_4539:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(39));
	CUT_4540:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(40));
	CUT_4541:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(41));
	CUT_4542:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(42));
	CUT_4543:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(43));
	CUT_4544:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(44));
	CUT_4545:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(45));
	CUT_4546:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(46));
	CUT_4547:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(47));
	CUT_4548:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(48));
	CUT_4549:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(90)(49));
	CUT_4550:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(0));
	CUT_4551:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(1));
	CUT_4552:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(2));
	CUT_4553:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(3));
	CUT_4554:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(4));
	CUT_4555:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(5));
	CUT_4556:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(6));
	CUT_4557:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(7));
	CUT_4558:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(8));
	CUT_4559:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(9));
	CUT_4560:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(10));
	CUT_4561:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(11));
	CUT_4562:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(12));
	CUT_4563:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(13));
	CUT_4564:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(14));
	CUT_4565:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(15));
	CUT_4566:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(16));
	CUT_4567:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(17));
	CUT_4568:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(18));
	CUT_4569:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(19));
	CUT_4570:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(20));
	CUT_4571:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(21));
	CUT_4572:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(22));
	CUT_4573:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(23));
	CUT_4574:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(24));
	CUT_4575:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(25));
	CUT_4576:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(26));
	CUT_4577:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(27));
	CUT_4578:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(28));
	CUT_4579:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(29));
	CUT_4580:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(30));
	CUT_4581:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(31));
	CUT_4582:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(32));
	CUT_4583:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(33));
	CUT_4584:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(34));
	CUT_4585:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(35));
	CUT_4586:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(36));
	CUT_4587:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(37));
	CUT_4588:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(38));
	CUT_4589:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(39));
	CUT_4590:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(40));
	CUT_4591:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(41));
	CUT_4592:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(42));
	CUT_4593:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(43));
	CUT_4594:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(44));
	CUT_4595:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(45));
	CUT_4596:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(46));
	CUT_4597:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(47));
	CUT_4598:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(48));
	CUT_4599:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(91)(49));
	CUT_4600:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(0));
	CUT_4601:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(1));
	CUT_4602:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(2));
	CUT_4603:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(3));
	CUT_4604:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(4));
	CUT_4605:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(5));
	CUT_4606:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(6));
	CUT_4607:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(7));
	CUT_4608:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(8));
	CUT_4609:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(9));
	CUT_4610:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(10));
	CUT_4611:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(11));
	CUT_4612:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(12));
	CUT_4613:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(13));
	CUT_4614:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(14));
	CUT_4615:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(15));
	CUT_4616:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(16));
	CUT_4617:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(17));
	CUT_4618:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(18));
	CUT_4619:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(19));
	CUT_4620:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(20));
	CUT_4621:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(21));
	CUT_4622:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(22));
	CUT_4623:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(23));
	CUT_4624:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(24));
	CUT_4625:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(25));
	CUT_4626:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(26));
	CUT_4627:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(27));
	CUT_4628:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(28));
	CUT_4629:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(29));
	CUT_4630:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(30));
	CUT_4631:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(31));
	CUT_4632:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(32));
	CUT_4633:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(33));
	CUT_4634:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(34));
	CUT_4635:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(35));
	CUT_4636:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(36));
	CUT_4637:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(37));
	CUT_4638:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(38));
	CUT_4639:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(39));
	CUT_4640:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(40));
	CUT_4641:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(41));
	CUT_4642:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(42));
	CUT_4643:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(43));
	CUT_4644:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(44));
	CUT_4645:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(45));
	CUT_4646:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(46));
	CUT_4647:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(47));
	CUT_4648:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(48));
	CUT_4649:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(92)(49));
	CUT_4650:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(0));
	CUT_4651:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(1));
	CUT_4652:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(2));
	CUT_4653:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(3));
	CUT_4654:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(4));
	CUT_4655:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(5));
	CUT_4656:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(6));
	CUT_4657:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(7));
	CUT_4658:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(8));
	CUT_4659:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(9));
	CUT_4660:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(10));
	CUT_4661:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(11));
	CUT_4662:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(12));
	CUT_4663:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(13));
	CUT_4664:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(14));
	CUT_4665:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(15));
	CUT_4666:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(16));
	CUT_4667:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(17));
	CUT_4668:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(18));
	CUT_4669:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(19));
	CUT_4670:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(20));
	CUT_4671:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(21));
	CUT_4672:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(22));
	CUT_4673:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(23));
	CUT_4674:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(24));
	CUT_4675:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(25));
	CUT_4676:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(26));
	CUT_4677:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(27));
	CUT_4678:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(28));
	CUT_4679:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(29));
	CUT_4680:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(30));
	CUT_4681:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(31));
	CUT_4682:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(32));
	CUT_4683:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(33));
	CUT_4684:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(34));
	CUT_4685:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(35));
	CUT_4686:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(36));
	CUT_4687:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(37));
	CUT_4688:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(38));
	CUT_4689:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(39));
	CUT_4690:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(40));
	CUT_4691:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(41));
	CUT_4692:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(42));
	CUT_4693:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(43));
	CUT_4694:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(44));
	CUT_4695:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(45));
	CUT_4696:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(46));
	CUT_4697:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(47));
	CUT_4698:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(48));
	CUT_4699:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(93)(49));
	CUT_4700:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(0));
	CUT_4701:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(1));
	CUT_4702:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(2));
	CUT_4703:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(3));
	CUT_4704:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(4));
	CUT_4705:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(5));
	CUT_4706:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(6));
	CUT_4707:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(7));
	CUT_4708:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(8));
	CUT_4709:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(9));
	CUT_4710:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(10));
	CUT_4711:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(11));
	CUT_4712:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(12));
	CUT_4713:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(13));
	CUT_4714:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(14));
	CUT_4715:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(15));
	CUT_4716:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(16));
	CUT_4717:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(17));
	CUT_4718:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(18));
	CUT_4719:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(19));
	CUT_4720:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(20));
	CUT_4721:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(21));
	CUT_4722:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(22));
	CUT_4723:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(23));
	CUT_4724:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(24));
	CUT_4725:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(25));
	CUT_4726:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(26));
	CUT_4727:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(27));
	CUT_4728:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(28));
	CUT_4729:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(29));
	CUT_4730:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(30));
	CUT_4731:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(31));
	CUT_4732:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(32));
	CUT_4733:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(33));
	CUT_4734:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(34));
	CUT_4735:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(35));
	CUT_4736:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(36));
	CUT_4737:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(37));
	CUT_4738:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(38));
	CUT_4739:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(39));
	CUT_4740:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(40));
	CUT_4741:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(41));
	CUT_4742:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(42));
	CUT_4743:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(43));
	CUT_4744:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(44));
	CUT_4745:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(45));
	CUT_4746:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(46));
	CUT_4747:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(47));
	CUT_4748:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(48));
	CUT_4749:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(94)(49));
	CUT_4750:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(0));
	CUT_4751:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(1));
	CUT_4752:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(2));
	CUT_4753:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(3));
	CUT_4754:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(4));
	CUT_4755:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(5));
	CUT_4756:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(6));
	CUT_4757:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(7));
	CUT_4758:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(8));
	CUT_4759:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(9));
	CUT_4760:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(10));
	CUT_4761:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(11));
	CUT_4762:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(12));
	CUT_4763:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(13));
	CUT_4764:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(14));
	CUT_4765:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(15));
	CUT_4766:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(16));
	CUT_4767:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(17));
	CUT_4768:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(18));
	CUT_4769:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(19));
	CUT_4770:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(20));
	CUT_4771:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(21));
	CUT_4772:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(22));
	CUT_4773:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(23));
	CUT_4774:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(24));
	CUT_4775:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(25));
	CUT_4776:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(26));
	CUT_4777:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(27));
	CUT_4778:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(28));
	CUT_4779:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(29));
	CUT_4780:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(30));
	CUT_4781:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(31));
	CUT_4782:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(32));
	CUT_4783:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(33));
	CUT_4784:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(34));
	CUT_4785:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(35));
	CUT_4786:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(36));
	CUT_4787:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(37));
	CUT_4788:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(38));
	CUT_4789:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(39));
	CUT_4790:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(40));
	CUT_4791:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(41));
	CUT_4792:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(42));
	CUT_4793:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(43));
	CUT_4794:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(44));
	CUT_4795:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(45));
	CUT_4796:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(46));
	CUT_4797:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(47));
	CUT_4798:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(48));
	CUT_4799:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(95)(49));
	CUT_4800:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(0));
	CUT_4801:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(1));
	CUT_4802:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(2));
	CUT_4803:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(3));
	CUT_4804:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(4));
	CUT_4805:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(5));
	CUT_4806:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(6));
	CUT_4807:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(7));
	CUT_4808:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(8));
	CUT_4809:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(9));
	CUT_4810:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(10));
	CUT_4811:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(11));
	CUT_4812:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(12));
	CUT_4813:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(13));
	CUT_4814:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(14));
	CUT_4815:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(15));
	CUT_4816:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(16));
	CUT_4817:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(17));
	CUT_4818:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(18));
	CUT_4819:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(19));
	CUT_4820:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(20));
	CUT_4821:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(21));
	CUT_4822:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(22));
	CUT_4823:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(23));
	CUT_4824:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(24));
	CUT_4825:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(25));
	CUT_4826:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(26));
	CUT_4827:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(27));
	CUT_4828:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(28));
	CUT_4829:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(29));
	CUT_4830:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(30));
	CUT_4831:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(31));
	CUT_4832:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(32));
	CUT_4833:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(33));
	CUT_4834:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(34));
	CUT_4835:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(35));
	CUT_4836:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(36));
	CUT_4837:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(37));
	CUT_4838:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(38));
	CUT_4839:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(39));
	CUT_4840:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(40));
	CUT_4841:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(41));
	CUT_4842:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(42));
	CUT_4843:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(43));
	CUT_4844:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(44));
	CUT_4845:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(45));
	CUT_4846:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(46));
	CUT_4847:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(47));
	CUT_4848:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(48));
	CUT_4849:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(96)(49));
	CUT_4850:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(0));
	CUT_4851:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(1));
	CUT_4852:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(2));
	CUT_4853:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(3));
	CUT_4854:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(4));
	CUT_4855:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(5));
	CUT_4856:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(6));
	CUT_4857:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(7));
	CUT_4858:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(8));
	CUT_4859:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(9));
	CUT_4860:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(10));
	CUT_4861:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(11));
	CUT_4862:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(12));
	CUT_4863:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(13));
	CUT_4864:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(14));
	CUT_4865:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(15));
	CUT_4866:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(16));
	CUT_4867:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(17));
	CUT_4868:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(18));
	CUT_4869:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(19));
	CUT_4870:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(20));
	CUT_4871:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(21));
	CUT_4872:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(22));
	CUT_4873:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(23));
	CUT_4874:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(24));
	CUT_4875:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(25));
	CUT_4876:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(26));
	CUT_4877:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(27));
	CUT_4878:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(28));
	CUT_4879:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(29));
	CUT_4880:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(30));
	CUT_4881:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(31));
	CUT_4882:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(32));
	CUT_4883:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(33));
	CUT_4884:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(34));
	CUT_4885:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(35));
	CUT_4886:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(36));
	CUT_4887:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(37));
	CUT_4888:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(38));
	CUT_4889:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(39));
	CUT_4890:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(40));
	CUT_4891:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(41));
	CUT_4892:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(42));
	CUT_4893:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(43));
	CUT_4894:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(44));
	CUT_4895:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(45));
	CUT_4896:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(46));
	CUT_4897:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(47));
	CUT_4898:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(48));
	CUT_4899:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(97)(49));
	CUT_4900:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(0));
	CUT_4901:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(1));
	CUT_4902:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(2));
	CUT_4903:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(3));
	CUT_4904:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(4));
	CUT_4905:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(5));
	CUT_4906:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(6));
	CUT_4907:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(7));
	CUT_4908:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(8));
	CUT_4909:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(9));
	CUT_4910:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(10));
	CUT_4911:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(11));
	CUT_4912:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(12));
	CUT_4913:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(13));
	CUT_4914:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(14));
	CUT_4915:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(15));
	CUT_4916:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(16));
	CUT_4917:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(17));
	CUT_4918:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(18));
	CUT_4919:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(19));
	CUT_4920:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(20));
	CUT_4921:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(21));
	CUT_4922:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(22));
	CUT_4923:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(23));
	CUT_4924:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(24));
	CUT_4925:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(25));
	CUT_4926:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(26));
	CUT_4927:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(27));
	CUT_4928:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(28));
	CUT_4929:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(29));
	CUT_4930:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(30));
	CUT_4931:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(31));
	CUT_4932:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(32));
	CUT_4933:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(33));
	CUT_4934:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(34));
	CUT_4935:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(35));
	CUT_4936:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(36));
	CUT_4937:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(37));
	CUT_4938:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(38));
	CUT_4939:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(39));
	CUT_4940:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(40));
	CUT_4941:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(41));
	CUT_4942:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(42));
	CUT_4943:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(43));
	CUT_4944:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(44));
	CUT_4945:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(45));
	CUT_4946:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(46));
	CUT_4947:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(47));
	CUT_4948:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(48));
	CUT_4949:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(98)(49));
	CUT_4950:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(0));
	CUT_4951:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(1));
	CUT_4952:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(2));
	CUT_4953:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(3));
	CUT_4954:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(4));
	CUT_4955:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(5));
	CUT_4956:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(6));
	CUT_4957:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(7));
	CUT_4958:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(8));
	CUT_4959:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(9));
	CUT_4960:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(10));
	CUT_4961:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(11));
	CUT_4962:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(12));
	CUT_4963:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(13));
	CUT_4964:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(14));
	CUT_4965:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(15));
	CUT_4966:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(16));
	CUT_4967:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(17));
	CUT_4968:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(18));
	CUT_4969:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(19));
	CUT_4970:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(20));
	CUT_4971:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(21));
	CUT_4972:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(22));
	CUT_4973:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(23));
	CUT_4974:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(24));
	CUT_4975:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(25));
	CUT_4976:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(26));
	CUT_4977:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(27));
	CUT_4978:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(28));
	CUT_4979:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(29));
	CUT_4980:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(30));
	CUT_4981:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(31));
	CUT_4982:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(32));
	CUT_4983:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(33));
	CUT_4984:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(34));
	CUT_4985:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(35));
	CUT_4986:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(36));
	CUT_4987:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(37));
	CUT_4988:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(38));
	CUT_4989:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(39));
	CUT_4990:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(40));
	CUT_4991:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(41));
	CUT_4992:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(42));
	CUT_4993:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(43));
	CUT_4994:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(44));
	CUT_4995:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(45));
	CUT_4996:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(46));
	CUT_4997:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(47));
	CUT_4998:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(48));
	CUT_4999:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(99)(49));
	CUT_5000:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(0));
	CUT_5001:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(1));
	CUT_5002:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(2));
	CUT_5003:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(3));
	CUT_5004:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(4));
	CUT_5005:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(5));
	CUT_5006:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(6));
	CUT_5007:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(7));
	CUT_5008:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(8));
	CUT_5009:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(9));
	CUT_5010:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(10));
	CUT_5011:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(11));
	CUT_5012:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(12));
	CUT_5013:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(13));
	CUT_5014:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(14));
	CUT_5015:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(15));
	CUT_5016:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(16));
	CUT_5017:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(17));
	CUT_5018:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(18));
	CUT_5019:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(19));
	CUT_5020:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(20));
	CUT_5021:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(21));
	CUT_5022:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(22));
	CUT_5023:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(23));
	CUT_5024:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(24));
	CUT_5025:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(25));
	CUT_5026:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(26));
	CUT_5027:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(27));
	CUT_5028:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(28));
	CUT_5029:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(29));
	CUT_5030:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(30));
	CUT_5031:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(31));
	CUT_5032:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(32));
	CUT_5033:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(33));
	CUT_5034:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(34));
	CUT_5035:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(35));
	CUT_5036:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(36));
	CUT_5037:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(37));
	CUT_5038:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(38));
	CUT_5039:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(39));
	CUT_5040:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(40));
	CUT_5041:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(41));
	CUT_5042:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(42));
	CUT_5043:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(43));
	CUT_5044:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(44));
	CUT_5045:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(45));
	CUT_5046:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(46));
	CUT_5047:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(47));
	CUT_5048:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(48));
	CUT_5049:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(100)(49));
	CUT_5050:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(0));
	CUT_5051:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(1));
	CUT_5052:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(2));
	CUT_5053:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(3));
	CUT_5054:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(4));
	CUT_5055:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(5));
	CUT_5056:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(6));
	CUT_5057:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(7));
	CUT_5058:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(8));
	CUT_5059:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(9));
	CUT_5060:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(10));
	CUT_5061:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(11));
	CUT_5062:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(12));
	CUT_5063:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(13));
	CUT_5064:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(14));
	CUT_5065:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(15));
	CUT_5066:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(16));
	CUT_5067:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(17));
	CUT_5068:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(18));
	CUT_5069:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(19));
	CUT_5070:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(20));
	CUT_5071:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(21));
	CUT_5072:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(22));
	CUT_5073:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(23));
	CUT_5074:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(24));
	CUT_5075:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(25));
	CUT_5076:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(26));
	CUT_5077:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(27));
	CUT_5078:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(28));
	CUT_5079:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(29));
	CUT_5080:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(30));
	CUT_5081:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(31));
	CUT_5082:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(32));
	CUT_5083:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(33));
	CUT_5084:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(34));
	CUT_5085:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(35));
	CUT_5086:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(36));
	CUT_5087:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(37));
	CUT_5088:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(38));
	CUT_5089:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(39));
	CUT_5090:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(40));
	CUT_5091:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(41));
	CUT_5092:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(42));
	CUT_5093:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(43));
	CUT_5094:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(44));
	CUT_5095:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(45));
	CUT_5096:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(46));
	CUT_5097:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(47));
	CUT_5098:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(48));
	CUT_5099:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(101)(49));
	CUT_5100:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(0));
	CUT_5101:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(1));
	CUT_5102:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(2));
	CUT_5103:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(3));
	CUT_5104:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(4));
	CUT_5105:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(5));
	CUT_5106:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(6));
	CUT_5107:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(7));
	CUT_5108:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(8));
	CUT_5109:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(9));
	CUT_5110:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(10));
	CUT_5111:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(11));
	CUT_5112:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(12));
	CUT_5113:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(13));
	CUT_5114:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(14));
	CUT_5115:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(15));
	CUT_5116:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(16));
	CUT_5117:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(17));
	CUT_5118:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(18));
	CUT_5119:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(19));
	CUT_5120:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(20));
	CUT_5121:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(21));
	CUT_5122:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(22));
	CUT_5123:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(23));
	CUT_5124:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(24));
	CUT_5125:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(25));
	CUT_5126:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(26));
	CUT_5127:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(27));
	CUT_5128:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(28));
	CUT_5129:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(29));
	CUT_5130:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(30));
	CUT_5131:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(31));
	CUT_5132:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(32));
	CUT_5133:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(33));
	CUT_5134:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(34));
	CUT_5135:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(35));
	CUT_5136:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(36));
	CUT_5137:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(37));
	CUT_5138:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(38));
	CUT_5139:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(39));
	CUT_5140:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(40));
	CUT_5141:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(41));
	CUT_5142:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(42));
	CUT_5143:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(43));
	CUT_5144:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(44));
	CUT_5145:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(45));
	CUT_5146:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(46));
	CUT_5147:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(47));
	CUT_5148:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(48));
	CUT_5149:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(102)(49));
	CUT_5150:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(0));
	CUT_5151:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(1));
	CUT_5152:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(2));
	CUT_5153:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(3));
	CUT_5154:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(4));
	CUT_5155:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(5));
	CUT_5156:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(6));
	CUT_5157:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(7));
	CUT_5158:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(8));
	CUT_5159:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(9));
	CUT_5160:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(10));
	CUT_5161:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(11));
	CUT_5162:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(12));
	CUT_5163:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(13));
	CUT_5164:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(14));
	CUT_5165:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(15));
	CUT_5166:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(16));
	CUT_5167:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(17));
	CUT_5168:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(18));
	CUT_5169:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(19));
	CUT_5170:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(20));
	CUT_5171:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(21));
	CUT_5172:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(22));
	CUT_5173:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(23));
	CUT_5174:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(24));
	CUT_5175:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(25));
	CUT_5176:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(26));
	CUT_5177:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(27));
	CUT_5178:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(28));
	CUT_5179:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(29));
	CUT_5180:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(30));
	CUT_5181:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(31));
	CUT_5182:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(32));
	CUT_5183:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(33));
	CUT_5184:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(34));
	CUT_5185:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(35));
	CUT_5186:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(36));
	CUT_5187:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(37));
	CUT_5188:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(38));
	CUT_5189:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(39));
	CUT_5190:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(40));
	CUT_5191:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(41));
	CUT_5192:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(42));
	CUT_5193:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(43));
	CUT_5194:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(44));
	CUT_5195:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(45));
	CUT_5196:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(46));
	CUT_5197:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(47));
	CUT_5198:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(48));
	CUT_5199:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(103)(49));
	CUT_5200:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(0));
	CUT_5201:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(1));
	CUT_5202:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(2));
	CUT_5203:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(3));
	CUT_5204:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(4));
	CUT_5205:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(5));
	CUT_5206:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(6));
	CUT_5207:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(7));
	CUT_5208:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(8));
	CUT_5209:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(9));
	CUT_5210:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(10));
	CUT_5211:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(11));
	CUT_5212:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(12));
	CUT_5213:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(13));
	CUT_5214:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(14));
	CUT_5215:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(15));
	CUT_5216:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(16));
	CUT_5217:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(17));
	CUT_5218:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(18));
	CUT_5219:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(19));
	CUT_5220:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(20));
	CUT_5221:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(21));
	CUT_5222:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(22));
	CUT_5223:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(23));
	CUT_5224:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(24));
	CUT_5225:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(25));
	CUT_5226:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(26));
	CUT_5227:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(27));
	CUT_5228:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(28));
	CUT_5229:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(29));
	CUT_5230:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(30));
	CUT_5231:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(31));
	CUT_5232:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(32));
	CUT_5233:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(33));
	CUT_5234:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(34));
	CUT_5235:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(35));
	CUT_5236:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(36));
	CUT_5237:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(37));
	CUT_5238:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(38));
	CUT_5239:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(39));
	CUT_5240:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(40));
	CUT_5241:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(41));
	CUT_5242:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(42));
	CUT_5243:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(43));
	CUT_5244:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(44));
	CUT_5245:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(45));
	CUT_5246:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(46));
	CUT_5247:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(47));
	CUT_5248:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(48));
	CUT_5249:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(104)(49));
	CUT_5250:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(0));
	CUT_5251:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(1));
	CUT_5252:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(2));
	CUT_5253:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(3));
	CUT_5254:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(4));
	CUT_5255:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(5));
	CUT_5256:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(6));
	CUT_5257:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(7));
	CUT_5258:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(8));
	CUT_5259:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(9));
	CUT_5260:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(10));
	CUT_5261:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(11));
	CUT_5262:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(12));
	CUT_5263:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(13));
	CUT_5264:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(14));
	CUT_5265:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(15));
	CUT_5266:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(16));
	CUT_5267:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(17));
	CUT_5268:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(18));
	CUT_5269:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(19));
	CUT_5270:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(20));
	CUT_5271:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(21));
	CUT_5272:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(22));
	CUT_5273:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(23));
	CUT_5274:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(24));
	CUT_5275:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(25));
	CUT_5276:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(26));
	CUT_5277:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(27));
	CUT_5278:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(28));
	CUT_5279:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(29));
	CUT_5280:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(30));
	CUT_5281:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(31));
	CUT_5282:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(32));
	CUT_5283:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(33));
	CUT_5284:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(34));
	CUT_5285:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(35));
	CUT_5286:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(36));
	CUT_5287:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(37));
	CUT_5288:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(38));
	CUT_5289:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(39));
	CUT_5290:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(40));
	CUT_5291:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(41));
	CUT_5292:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(42));
	CUT_5293:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(43));
	CUT_5294:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(44));
	CUT_5295:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(45));
	CUT_5296:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(46));
	CUT_5297:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(47));
	CUT_5298:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(48));
	CUT_5299:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(105)(49));
	CUT_5300:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(0));
	CUT_5301:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(1));
	CUT_5302:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(2));
	CUT_5303:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(3));
	CUT_5304:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(4));
	CUT_5305:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(5));
	CUT_5306:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(6));
	CUT_5307:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(7));
	CUT_5308:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(8));
	CUT_5309:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(9));
	CUT_5310:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(10));
	CUT_5311:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(11));
	CUT_5312:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(12));
	CUT_5313:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(13));
	CUT_5314:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(14));
	CUT_5315:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(15));
	CUT_5316:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(16));
	CUT_5317:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(17));
	CUT_5318:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(18));
	CUT_5319:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(19));
	CUT_5320:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(20));
	CUT_5321:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(21));
	CUT_5322:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(22));
	CUT_5323:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(23));
	CUT_5324:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(24));
	CUT_5325:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(25));
	CUT_5326:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(26));
	CUT_5327:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(27));
	CUT_5328:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(28));
	CUT_5329:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(29));
	CUT_5330:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(30));
	CUT_5331:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(31));
	CUT_5332:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(32));
	CUT_5333:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(33));
	CUT_5334:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(34));
	CUT_5335:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(35));
	CUT_5336:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(36));
	CUT_5337:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(37));
	CUT_5338:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(38));
	CUT_5339:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(39));
	CUT_5340:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(40));
	CUT_5341:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(41));
	CUT_5342:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(42));
	CUT_5343:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(43));
	CUT_5344:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(44));
	CUT_5345:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(45));
	CUT_5346:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(46));
	CUT_5347:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(47));
	CUT_5348:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(48));
	CUT_5349:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(106)(49));
	CUT_5350:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(0));
	CUT_5351:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(1));
	CUT_5352:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(2));
	CUT_5353:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(3));
	CUT_5354:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(4));
	CUT_5355:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(5));
	CUT_5356:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(6));
	CUT_5357:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(7));
	CUT_5358:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(8));
	CUT_5359:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(9));
	CUT_5360:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(10));
	CUT_5361:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(11));
	CUT_5362:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(12));
	CUT_5363:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(13));
	CUT_5364:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(14));
	CUT_5365:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(15));
	CUT_5366:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(16));
	CUT_5367:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(17));
	CUT_5368:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(18));
	CUT_5369:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(19));
	CUT_5370:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(20));
	CUT_5371:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(21));
	CUT_5372:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(22));
	CUT_5373:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(23));
	CUT_5374:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(24));
	CUT_5375:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(25));
	CUT_5376:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(26));
	CUT_5377:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(27));
	CUT_5378:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(28));
	CUT_5379:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(29));
	CUT_5380:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(30));
	CUT_5381:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(31));
	CUT_5382:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(32));
	CUT_5383:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(33));
	CUT_5384:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(34));
	CUT_5385:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(35));
	CUT_5386:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(36));
	CUT_5387:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(37));
	CUT_5388:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(38));
	CUT_5389:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(39));
	CUT_5390:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(40));
	CUT_5391:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(41));
	CUT_5392:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(42));
	CUT_5393:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(43));
	CUT_5394:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(44));
	CUT_5395:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(45));
	CUT_5396:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(46));
	CUT_5397:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(47));
	CUT_5398:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(48));
	CUT_5399:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(107)(49));
	CUT_5400:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(0));
	CUT_5401:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(1));
	CUT_5402:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(2));
	CUT_5403:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(3));
	CUT_5404:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(4));
	CUT_5405:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(5));
	CUT_5406:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(6));
	CUT_5407:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(7));
	CUT_5408:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(8));
	CUT_5409:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(9));
	CUT_5410:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(10));
	CUT_5411:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(11));
	CUT_5412:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(12));
	CUT_5413:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(13));
	CUT_5414:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(14));
	CUT_5415:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(15));
	CUT_5416:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(16));
	CUT_5417:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(17));
	CUT_5418:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(18));
	CUT_5419:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(19));
	CUT_5420:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(20));
	CUT_5421:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(21));
	CUT_5422:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(22));
	CUT_5423:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(23));
	CUT_5424:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(24));
	CUT_5425:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(25));
	CUT_5426:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(26));
	CUT_5427:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(27));
	CUT_5428:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(28));
	CUT_5429:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(29));
	CUT_5430:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(30));
	CUT_5431:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(31));
	CUT_5432:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(32));
	CUT_5433:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(33));
	CUT_5434:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(34));
	CUT_5435:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(35));
	CUT_5436:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(36));
	CUT_5437:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(37));
	CUT_5438:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(38));
	CUT_5439:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(39));
	CUT_5440:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(40));
	CUT_5441:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(41));
	CUT_5442:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(42));
	CUT_5443:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(43));
	CUT_5444:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(44));
	CUT_5445:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(45));
	CUT_5446:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(46));
	CUT_5447:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(47));
	CUT_5448:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(48));
	CUT_5449:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(108)(49));
	CUT_5450:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(0));
	CUT_5451:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(1));
	CUT_5452:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(2));
	CUT_5453:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(3));
	CUT_5454:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(4));
	CUT_5455:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(5));
	CUT_5456:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(6));
	CUT_5457:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(7));
	CUT_5458:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(8));
	CUT_5459:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(9));
	CUT_5460:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(10));
	CUT_5461:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(11));
	CUT_5462:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(12));
	CUT_5463:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(13));
	CUT_5464:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(14));
	CUT_5465:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(15));
	CUT_5466:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(16));
	CUT_5467:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(17));
	CUT_5468:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(18));
	CUT_5469:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(19));
	CUT_5470:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(20));
	CUT_5471:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(21));
	CUT_5472:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(22));
	CUT_5473:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(23));
	CUT_5474:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(24));
	CUT_5475:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(25));
	CUT_5476:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(26));
	CUT_5477:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(27));
	CUT_5478:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(28));
	CUT_5479:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(29));
	CUT_5480:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(30));
	CUT_5481:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(31));
	CUT_5482:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(32));
	CUT_5483:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(33));
	CUT_5484:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(34));
	CUT_5485:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(35));
	CUT_5486:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(36));
	CUT_5487:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(37));
	CUT_5488:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(38));
	CUT_5489:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(39));
	CUT_5490:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(40));
	CUT_5491:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(41));
	CUT_5492:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(42));
	CUT_5493:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(43));
	CUT_5494:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(44));
	CUT_5495:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(45));
	CUT_5496:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(46));
	CUT_5497:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(47));
	CUT_5498:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(48));
	CUT_5499:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(109)(49));
	CUT_5500:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(0));
	CUT_5501:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(1));
	CUT_5502:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(2));
	CUT_5503:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(3));
	CUT_5504:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(4));
	CUT_5505:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(5));
	CUT_5506:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(6));
	CUT_5507:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(7));
	CUT_5508:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(8));
	CUT_5509:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(9));
	CUT_5510:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(10));
	CUT_5511:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(11));
	CUT_5512:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(12));
	CUT_5513:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(13));
	CUT_5514:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(14));
	CUT_5515:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(15));
	CUT_5516:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(16));
	CUT_5517:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(17));
	CUT_5518:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(18));
	CUT_5519:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(19));
	CUT_5520:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(20));
	CUT_5521:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(21));
	CUT_5522:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(22));
	CUT_5523:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(23));
	CUT_5524:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(24));
	CUT_5525:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(25));
	CUT_5526:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(26));
	CUT_5527:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(27));
	CUT_5528:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(28));
	CUT_5529:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(29));
	CUT_5530:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(30));
	CUT_5531:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(31));
	CUT_5532:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(32));
	CUT_5533:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(33));
	CUT_5534:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(34));
	CUT_5535:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(35));
	CUT_5536:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(36));
	CUT_5537:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(37));
	CUT_5538:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(38));
	CUT_5539:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(39));
	CUT_5540:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(40));
	CUT_5541:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(41));
	CUT_5542:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(42));
	CUT_5543:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(43));
	CUT_5544:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(44));
	CUT_5545:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(45));
	CUT_5546:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(46));
	CUT_5547:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(47));
	CUT_5548:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(48));
	CUT_5549:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(110)(49));
	CUT_5550:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(0));
	CUT_5551:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(1));
	CUT_5552:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(2));
	CUT_5553:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(3));
	CUT_5554:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(4));
	CUT_5555:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(5));
	CUT_5556:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(6));
	CUT_5557:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(7));
	CUT_5558:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(8));
	CUT_5559:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(9));
	CUT_5560:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(10));
	CUT_5561:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(11));
	CUT_5562:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(12));
	CUT_5563:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(13));
	CUT_5564:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(14));
	CUT_5565:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(15));
	CUT_5566:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(16));
	CUT_5567:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(17));
	CUT_5568:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(18));
	CUT_5569:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(19));
	CUT_5570:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(20));
	CUT_5571:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(21));
	CUT_5572:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(22));
	CUT_5573:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(23));
	CUT_5574:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(24));
	CUT_5575:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(25));
	CUT_5576:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(26));
	CUT_5577:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(27));
	CUT_5578:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(28));
	CUT_5579:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(29));
	CUT_5580:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(30));
	CUT_5581:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(31));
	CUT_5582:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(32));
	CUT_5583:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(33));
	CUT_5584:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(34));
	CUT_5585:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(35));
	CUT_5586:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(36));
	CUT_5587:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(37));
	CUT_5588:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(38));
	CUT_5589:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(39));
	CUT_5590:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(40));
	CUT_5591:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(41));
	CUT_5592:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(42));
	CUT_5593:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(43));
	CUT_5594:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(44));
	CUT_5595:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(45));
	CUT_5596:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(46));
	CUT_5597:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(47));
	CUT_5598:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(48));
	CUT_5599:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(111)(49));
	CUT_5600:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(0));
	CUT_5601:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(1));
	CUT_5602:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(2));
	CUT_5603:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(3));
	CUT_5604:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(4));
	CUT_5605:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(5));
	CUT_5606:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(6));
	CUT_5607:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(7));
	CUT_5608:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(8));
	CUT_5609:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(9));
	CUT_5610:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(10));
	CUT_5611:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(11));
	CUT_5612:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(12));
	CUT_5613:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(13));
	CUT_5614:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(14));
	CUT_5615:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(15));
	CUT_5616:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(16));
	CUT_5617:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(17));
	CUT_5618:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(18));
	CUT_5619:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(19));
	CUT_5620:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(20));
	CUT_5621:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(21));
	CUT_5622:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(22));
	CUT_5623:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(23));
	CUT_5624:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(24));
	CUT_5625:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(25));
	CUT_5626:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(26));
	CUT_5627:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(27));
	CUT_5628:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(28));
	CUT_5629:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(29));
	CUT_5630:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(30));
	CUT_5631:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(31));
	CUT_5632:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(32));
	CUT_5633:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(33));
	CUT_5634:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(34));
	CUT_5635:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(35));
	CUT_5636:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(36));
	CUT_5637:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(37));
	CUT_5638:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(38));
	CUT_5639:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(39));
	CUT_5640:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(40));
	CUT_5641:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(41));
	CUT_5642:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(42));
	CUT_5643:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(43));
	CUT_5644:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(44));
	CUT_5645:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(45));
	CUT_5646:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(46));
	CUT_5647:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(47));
	CUT_5648:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(48));
	CUT_5649:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(112)(49));
	CUT_5650:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(0));
	CUT_5651:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(1));
	CUT_5652:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(2));
	CUT_5653:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(3));
	CUT_5654:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(4));
	CUT_5655:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(5));
	CUT_5656:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(6));
	CUT_5657:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(7));
	CUT_5658:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(8));
	CUT_5659:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(9));
	CUT_5660:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(10));
	CUT_5661:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(11));
	CUT_5662:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(12));
	CUT_5663:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(13));
	CUT_5664:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(14));
	CUT_5665:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(15));
	CUT_5666:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(16));
	CUT_5667:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(17));
	CUT_5668:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(18));
	CUT_5669:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(19));
	CUT_5670:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(20));
	CUT_5671:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(21));
	CUT_5672:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(22));
	CUT_5673:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(23));
	CUT_5674:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(24));
	CUT_5675:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(25));
	CUT_5676:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(26));
	CUT_5677:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(27));
	CUT_5678:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(28));
	CUT_5679:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(29));
	CUT_5680:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(30));
	CUT_5681:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(31));
	CUT_5682:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(32));
	CUT_5683:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(33));
	CUT_5684:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(34));
	CUT_5685:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(35));
	CUT_5686:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(36));
	CUT_5687:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(37));
	CUT_5688:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(38));
	CUT_5689:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(39));
	CUT_5690:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(40));
	CUT_5691:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(41));
	CUT_5692:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(42));
	CUT_5693:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(43));
	CUT_5694:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(44));
	CUT_5695:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(45));
	CUT_5696:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(46));
	CUT_5697:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(47));
	CUT_5698:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(48));
	CUT_5699:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(113)(49));
	CUT_5700:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(0));
	CUT_5701:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(1));
	CUT_5702:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(2));
	CUT_5703:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(3));
	CUT_5704:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(4));
	CUT_5705:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(5));
	CUT_5706:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(6));
	CUT_5707:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(7));
	CUT_5708:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(8));
	CUT_5709:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(9));
	CUT_5710:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(10));
	CUT_5711:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(11));
	CUT_5712:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(12));
	CUT_5713:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(13));
	CUT_5714:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(14));
	CUT_5715:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(15));
	CUT_5716:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(16));
	CUT_5717:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(17));
	CUT_5718:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(18));
	CUT_5719:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(19));
	CUT_5720:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(20));
	CUT_5721:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(21));
	CUT_5722:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(22));
	CUT_5723:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(23));
	CUT_5724:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(24));
	CUT_5725:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(25));
	CUT_5726:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(26));
	CUT_5727:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(27));
	CUT_5728:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(28));
	CUT_5729:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(29));
	CUT_5730:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(30));
	CUT_5731:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(31));
	CUT_5732:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(32));
	CUT_5733:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(33));
	CUT_5734:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(34));
	CUT_5735:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(35));
	CUT_5736:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(36));
	CUT_5737:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(37));
	CUT_5738:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(38));
	CUT_5739:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(39));
	CUT_5740:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(40));
	CUT_5741:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(41));
	CUT_5742:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(42));
	CUT_5743:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(43));
	CUT_5744:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(44));
	CUT_5745:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(45));
	CUT_5746:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(46));
	CUT_5747:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(47));
	CUT_5748:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(48));
	CUT_5749:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(114)(49));
	CUT_5750:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(0));
	CUT_5751:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(1));
	CUT_5752:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(2));
	CUT_5753:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(3));
	CUT_5754:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(4));
	CUT_5755:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(5));
	CUT_5756:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(6));
	CUT_5757:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(7));
	CUT_5758:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(8));
	CUT_5759:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(9));
	CUT_5760:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(10));
	CUT_5761:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(11));
	CUT_5762:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(12));
	CUT_5763:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(13));
	CUT_5764:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(14));
	CUT_5765:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(15));
	CUT_5766:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(16));
	CUT_5767:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(17));
	CUT_5768:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(18));
	CUT_5769:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(19));
	CUT_5770:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(20));
	CUT_5771:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(21));
	CUT_5772:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(22));
	CUT_5773:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(23));
	CUT_5774:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(24));
	CUT_5775:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(25));
	CUT_5776:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(26));
	CUT_5777:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(27));
	CUT_5778:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(28));
	CUT_5779:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(29));
	CUT_5780:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(30));
	CUT_5781:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(31));
	CUT_5782:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(32));
	CUT_5783:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(33));
	CUT_5784:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(34));
	CUT_5785:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(35));
	CUT_5786:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(36));
	CUT_5787:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(37));
	CUT_5788:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(38));
	CUT_5789:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(39));
	CUT_5790:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(40));
	CUT_5791:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(41));
	CUT_5792:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(42));
	CUT_5793:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(43));
	CUT_5794:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(44));
	CUT_5795:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(45));
	CUT_5796:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(46));
	CUT_5797:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(47));
	CUT_5798:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(48));
	CUT_5799:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(115)(49));
	CUT_5800:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(0));
	CUT_5801:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(1));
	CUT_5802:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(2));
	CUT_5803:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(3));
	CUT_5804:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(4));
	CUT_5805:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(5));
	CUT_5806:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(6));
	CUT_5807:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(7));
	CUT_5808:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(8));
	CUT_5809:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(9));
	CUT_5810:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(10));
	CUT_5811:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(11));
	CUT_5812:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(12));
	CUT_5813:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(13));
	CUT_5814:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(14));
	CUT_5815:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(15));
	CUT_5816:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(16));
	CUT_5817:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(17));
	CUT_5818:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(18));
	CUT_5819:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(19));
	CUT_5820:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(20));
	CUT_5821:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(21));
	CUT_5822:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(22));
	CUT_5823:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(23));
	CUT_5824:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(24));
	CUT_5825:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(25));
	CUT_5826:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(26));
	CUT_5827:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(27));
	CUT_5828:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(28));
	CUT_5829:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(29));
	CUT_5830:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(30));
	CUT_5831:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(31));
	CUT_5832:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(32));
	CUT_5833:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(33));
	CUT_5834:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(34));
	CUT_5835:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(35));
	CUT_5836:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(36));
	CUT_5837:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(37));
	CUT_5838:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(38));
	CUT_5839:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(39));
	CUT_5840:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(40));
	CUT_5841:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(41));
	CUT_5842:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(42));
	CUT_5843:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(43));
	CUT_5844:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(44));
	CUT_5845:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(45));
	CUT_5846:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(46));
	CUT_5847:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(47));
	CUT_5848:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(48));
	CUT_5849:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(116)(49));
	CUT_5850:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(0));
	CUT_5851:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(1));
	CUT_5852:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(2));
	CUT_5853:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(3));
	CUT_5854:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(4));
	CUT_5855:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(5));
	CUT_5856:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(6));
	CUT_5857:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(7));
	CUT_5858:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(8));
	CUT_5859:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(9));
	CUT_5860:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(10));
	CUT_5861:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(11));
	CUT_5862:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(12));
	CUT_5863:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(13));
	CUT_5864:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(14));
	CUT_5865:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(15));
	CUT_5866:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(16));
	CUT_5867:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(17));
	CUT_5868:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(18));
	CUT_5869:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(19));
	CUT_5870:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(20));
	CUT_5871:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(21));
	CUT_5872:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(22));
	CUT_5873:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(23));
	CUT_5874:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(24));
	CUT_5875:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(25));
	CUT_5876:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(26));
	CUT_5877:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(27));
	CUT_5878:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(28));
	CUT_5879:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(29));
	CUT_5880:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(30));
	CUT_5881:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(31));
	CUT_5882:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(32));
	CUT_5883:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(33));
	CUT_5884:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(34));
	CUT_5885:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(35));
	CUT_5886:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(36));
	CUT_5887:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(37));
	CUT_5888:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(38));
	CUT_5889:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(39));
	CUT_5890:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(40));
	CUT_5891:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(41));
	CUT_5892:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(42));
	CUT_5893:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(43));
	CUT_5894:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(44));
	CUT_5895:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(45));
	CUT_5896:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(46));
	CUT_5897:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(47));
	CUT_5898:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(48));
	CUT_5899:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(117)(49));
	CUT_5900:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(0));
	CUT_5901:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(1));
	CUT_5902:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(2));
	CUT_5903:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(3));
	CUT_5904:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(4));
	CUT_5905:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(5));
	CUT_5906:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(6));
	CUT_5907:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(7));
	CUT_5908:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(8));
	CUT_5909:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(9));
	CUT_5910:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(10));
	CUT_5911:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(11));
	CUT_5912:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(12));
	CUT_5913:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(13));
	CUT_5914:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(14));
	CUT_5915:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(15));
	CUT_5916:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(16));
	CUT_5917:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(17));
	CUT_5918:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(18));
	CUT_5919:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(19));
	CUT_5920:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(20));
	CUT_5921:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(21));
	CUT_5922:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(22));
	CUT_5923:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(23));
	CUT_5924:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(24));
	CUT_5925:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(25));
	CUT_5926:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(26));
	CUT_5927:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(27));
	CUT_5928:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(28));
	CUT_5929:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(29));
	CUT_5930:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(30));
	CUT_5931:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(31));
	CUT_5932:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(32));
	CUT_5933:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(33));
	CUT_5934:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(34));
	CUT_5935:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(35));
	CUT_5936:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(36));
	CUT_5937:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(37));
	CUT_5938:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(38));
	CUT_5939:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(39));
	CUT_5940:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(40));
	CUT_5941:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(41));
	CUT_5942:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(42));
	CUT_5943:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(43));
	CUT_5944:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(44));
	CUT_5945:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(45));
	CUT_5946:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(46));
	CUT_5947:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(47));
	CUT_5948:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(48));
	CUT_5949:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(118)(49));
	CUT_5950:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(0));
	CUT_5951:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(1));
	CUT_5952:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(2));
	CUT_5953:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(3));
	CUT_5954:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(4));
	CUT_5955:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(5));
	CUT_5956:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(6));
	CUT_5957:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(7));
	CUT_5958:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(8));
	CUT_5959:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(9));
	CUT_5960:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(10));
	CUT_5961:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(11));
	CUT_5962:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(12));
	CUT_5963:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(13));
	CUT_5964:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(14));
	CUT_5965:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(15));
	CUT_5966:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(16));
	CUT_5967:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(17));
	CUT_5968:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(18));
	CUT_5969:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(19));
	CUT_5970:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(20));
	CUT_5971:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(21));
	CUT_5972:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(22));
	CUT_5973:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(23));
	CUT_5974:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(24));
	CUT_5975:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(25));
	CUT_5976:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(26));
	CUT_5977:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(27));
	CUT_5978:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(28));
	CUT_5979:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(29));
	CUT_5980:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(30));
	CUT_5981:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(31));
	CUT_5982:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(32));
	CUT_5983:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(33));
	CUT_5984:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(34));
	CUT_5985:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(35));
	CUT_5986:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(36));
	CUT_5987:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(37));
	CUT_5988:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(38));
	CUT_5989:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(39));
	CUT_5990:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(40));
	CUT_5991:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(41));
	CUT_5992:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(42));
	CUT_5993:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(43));
	CUT_5994:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(44));
	CUT_5995:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(45));
	CUT_5996:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(46));
	CUT_5997:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(47));
	CUT_5998:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(48));
	CUT_5999:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(119)(49));
	CUT_6000:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(0));
	CUT_6001:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(1));
	CUT_6002:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(2));
	CUT_6003:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(3));
	CUT_6004:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(4));
	CUT_6005:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(5));
	CUT_6006:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(6));
	CUT_6007:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(7));
	CUT_6008:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(8));
	CUT_6009:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(9));
	CUT_6010:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(10));
	CUT_6011:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(11));
	CUT_6012:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(12));
	CUT_6013:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(13));
	CUT_6014:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(14));
	CUT_6015:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(15));
	CUT_6016:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(16));
	CUT_6017:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(17));
	CUT_6018:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(18));
	CUT_6019:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(19));
	CUT_6020:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(20));
	CUT_6021:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(21));
	CUT_6022:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(22));
	CUT_6023:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(23));
	CUT_6024:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(24));
	CUT_6025:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(25));
	CUT_6026:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(26));
	CUT_6027:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(27));
	CUT_6028:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(28));
	CUT_6029:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(29));
	CUT_6030:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(30));
	CUT_6031:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(31));
	CUT_6032:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(32));
	CUT_6033:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(33));
	CUT_6034:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(34));
	CUT_6035:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(35));
	CUT_6036:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(36));
	CUT_6037:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(37));
	CUT_6038:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(38));
	CUT_6039:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(39));
	CUT_6040:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(40));
	CUT_6041:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(41));
	CUT_6042:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(42));
	CUT_6043:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(43));
	CUT_6044:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(44));
	CUT_6045:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(45));
	CUT_6046:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(46));
	CUT_6047:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(47));
	CUT_6048:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(48));
	CUT_6049:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(120)(49));
	CUT_6050:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(0));
	CUT_6051:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(1));
	CUT_6052:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(2));
	CUT_6053:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(3));
	CUT_6054:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(4));
	CUT_6055:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(5));
	CUT_6056:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(6));
	CUT_6057:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(7));
	CUT_6058:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(8));
	CUT_6059:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(9));
	CUT_6060:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(10));
	CUT_6061:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(11));
	CUT_6062:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(12));
	CUT_6063:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(13));
	CUT_6064:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(14));
	CUT_6065:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(15));
	CUT_6066:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(16));
	CUT_6067:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(17));
	CUT_6068:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(18));
	CUT_6069:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(19));
	CUT_6070:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(20));
	CUT_6071:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(21));
	CUT_6072:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(22));
	CUT_6073:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(23));
	CUT_6074:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(24));
	CUT_6075:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(25));
	CUT_6076:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(26));
	CUT_6077:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(27));
	CUT_6078:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(28));
	CUT_6079:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(29));
	CUT_6080:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(30));
	CUT_6081:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(31));
	CUT_6082:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(32));
	CUT_6083:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(33));
	CUT_6084:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(34));
	CUT_6085:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(35));
	CUT_6086:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(36));
	CUT_6087:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(37));
	CUT_6088:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(38));
	CUT_6089:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(39));
	CUT_6090:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(40));
	CUT_6091:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(41));
	CUT_6092:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(42));
	CUT_6093:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(43));
	CUT_6094:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(44));
	CUT_6095:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(45));
	CUT_6096:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(46));
	CUT_6097:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(47));
	CUT_6098:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(48));
	CUT_6099:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(121)(49));
	CUT_6100:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(0));
	CUT_6101:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(1));
	CUT_6102:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(2));
	CUT_6103:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(3));
	CUT_6104:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(4));
	CUT_6105:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(5));
	CUT_6106:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(6));
	CUT_6107:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(7));
	CUT_6108:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(8));
	CUT_6109:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(9));
	CUT_6110:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(10));
	CUT_6111:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(11));
	CUT_6112:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(12));
	CUT_6113:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(13));
	CUT_6114:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(14));
	CUT_6115:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(15));
	CUT_6116:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(16));
	CUT_6117:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(17));
	CUT_6118:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(18));
	CUT_6119:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(19));
	CUT_6120:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(20));
	CUT_6121:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(21));
	CUT_6122:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(22));
	CUT_6123:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(23));
	CUT_6124:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(24));
	CUT_6125:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(25));
	CUT_6126:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(26));
	CUT_6127:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(27));
	CUT_6128:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(28));
	CUT_6129:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(29));
	CUT_6130:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(30));
	CUT_6131:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(31));
	CUT_6132:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(32));
	CUT_6133:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(33));
	CUT_6134:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(34));
	CUT_6135:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(35));
	CUT_6136:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(36));
	CUT_6137:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(37));
	CUT_6138:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(38));
	CUT_6139:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(39));
	CUT_6140:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(40));
	CUT_6141:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(41));
	CUT_6142:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(42));
	CUT_6143:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(43));
	CUT_6144:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(44));
	CUT_6145:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(45));
	CUT_6146:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(46));
	CUT_6147:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(47));
	CUT_6148:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(48));
	CUT_6149:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(122)(49));
	CUT_6150:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(0));
	CUT_6151:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(1));
	CUT_6152:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(2));
	CUT_6153:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(3));
	CUT_6154:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(4));
	CUT_6155:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(5));
	CUT_6156:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(6));
	CUT_6157:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(7));
	CUT_6158:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(8));
	CUT_6159:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(9));
	CUT_6160:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(10));
	CUT_6161:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(11));
	CUT_6162:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(12));
	CUT_6163:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(13));
	CUT_6164:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(14));
	CUT_6165:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(15));
	CUT_6166:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(16));
	CUT_6167:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(17));
	CUT_6168:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(18));
	CUT_6169:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(19));
	CUT_6170:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(20));
	CUT_6171:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(21));
	CUT_6172:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(22));
	CUT_6173:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(23));
	CUT_6174:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(24));
	CUT_6175:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(25));
	CUT_6176:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(26));
	CUT_6177:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(27));
	CUT_6178:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(28));
	CUT_6179:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(29));
	CUT_6180:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(30));
	CUT_6181:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(31));
	CUT_6182:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(32));
	CUT_6183:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(33));
	CUT_6184:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(34));
	CUT_6185:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(35));
	CUT_6186:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(36));
	CUT_6187:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(37));
	CUT_6188:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(38));
	CUT_6189:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(39));
	CUT_6190:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(40));
	CUT_6191:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(41));
	CUT_6192:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(42));
	CUT_6193:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(43));
	CUT_6194:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(44));
	CUT_6195:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(45));
	CUT_6196:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(46));
	CUT_6197:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(47));
	CUT_6198:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(48));
	CUT_6199:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(123)(49));
	CUT_6200:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(0));
	CUT_6201:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(1));
	CUT_6202:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(2));
	CUT_6203:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(3));
	CUT_6204:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(4));
	CUT_6205:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(5));
	CUT_6206:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(6));
	CUT_6207:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(7));
	CUT_6208:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(8));
	CUT_6209:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(9));
	CUT_6210:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(10));
	CUT_6211:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(11));
	CUT_6212:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(12));
	CUT_6213:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(13));
	CUT_6214:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(14));
	CUT_6215:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(15));
	CUT_6216:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(16));
	CUT_6217:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(17));
	CUT_6218:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(18));
	CUT_6219:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(19));
	CUT_6220:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(20));
	CUT_6221:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(21));
	CUT_6222:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(22));
	CUT_6223:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(23));
	CUT_6224:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(24));
	CUT_6225:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(25));
	CUT_6226:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(26));
	CUT_6227:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(27));
	CUT_6228:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(28));
	CUT_6229:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(29));
	CUT_6230:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(30));
	CUT_6231:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(31));
	CUT_6232:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(32));
	CUT_6233:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(33));
	CUT_6234:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(34));
	CUT_6235:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(35));
	CUT_6236:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(36));
	CUT_6237:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(37));
	CUT_6238:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(38));
	CUT_6239:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(39));
	CUT_6240:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(40));
	CUT_6241:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(41));
	CUT_6242:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(42));
	CUT_6243:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(43));
	CUT_6244:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(44));
	CUT_6245:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(45));
	CUT_6246:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(46));
	CUT_6247:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(47));
	CUT_6248:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(48));
	CUT_6249:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(124)(49));
	CUT_6250:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(0));
	CUT_6251:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(1));
	CUT_6252:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(2));
	CUT_6253:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(3));
	CUT_6254:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(4));
	CUT_6255:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(5));
	CUT_6256:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(6));
	CUT_6257:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(7));
	CUT_6258:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(8));
	CUT_6259:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(9));
	CUT_6260:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(10));
	CUT_6261:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(11));
	CUT_6262:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(12));
	CUT_6263:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(13));
	CUT_6264:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(14));
	CUT_6265:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(15));
	CUT_6266:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(16));
	CUT_6267:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(17));
	CUT_6268:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(18));
	CUT_6269:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(19));
	CUT_6270:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(20));
	CUT_6271:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(21));
	CUT_6272:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(22));
	CUT_6273:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(23));
	CUT_6274:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(24));
	CUT_6275:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(25));
	CUT_6276:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(26));
	CUT_6277:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(27));
	CUT_6278:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(28));
	CUT_6279:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(29));
	CUT_6280:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(30));
	CUT_6281:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(31));
	CUT_6282:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(32));
	CUT_6283:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(33));
	CUT_6284:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(34));
	CUT_6285:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(35));
	CUT_6286:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(36));
	CUT_6287:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(37));
	CUT_6288:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(38));
	CUT_6289:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(39));
	CUT_6290:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(40));
	CUT_6291:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(41));
	CUT_6292:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(42));
	CUT_6293:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(43));
	CUT_6294:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(44));
	CUT_6295:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(45));
	CUT_6296:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(46));
	CUT_6297:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(47));
	CUT_6298:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(48));
	CUT_6299:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(125)(49));
	CUT_6300:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(0));
	CUT_6301:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(1));
	CUT_6302:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(2));
	CUT_6303:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(3));
	CUT_6304:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(4));
	CUT_6305:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(5));
	CUT_6306:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(6));
	CUT_6307:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(7));
	CUT_6308:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(8));
	CUT_6309:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(9));
	CUT_6310:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(10));
	CUT_6311:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(11));
	CUT_6312:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(12));
	CUT_6313:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(13));
	CUT_6314:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(14));
	CUT_6315:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(15));
	CUT_6316:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(16));
	CUT_6317:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(17));
	CUT_6318:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(18));
	CUT_6319:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(19));
	CUT_6320:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(20));
	CUT_6321:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(21));
	CUT_6322:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(22));
	CUT_6323:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(23));
	CUT_6324:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(24));
	CUT_6325:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(25));
	CUT_6326:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(26));
	CUT_6327:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(27));
	CUT_6328:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(28));
	CUT_6329:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(29));
	CUT_6330:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(30));
	CUT_6331:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(31));
	CUT_6332:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(32));
	CUT_6333:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(33));
	CUT_6334:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(34));
	CUT_6335:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(35));
	CUT_6336:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(36));
	CUT_6337:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(37));
	CUT_6338:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(38));
	CUT_6339:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(39));
	CUT_6340:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(40));
	CUT_6341:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(41));
	CUT_6342:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(42));
	CUT_6343:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(43));
	CUT_6344:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(44));
	CUT_6345:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(45));
	CUT_6346:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(46));
	CUT_6347:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(47));
	CUT_6348:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(48));
	CUT_6349:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(126)(49));
	CUT_6350:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(0));
	CUT_6351:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(1));
	CUT_6352:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(2));
	CUT_6353:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(3));
	CUT_6354:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(4));
	CUT_6355:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(5));
	CUT_6356:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(6));
	CUT_6357:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(7));
	CUT_6358:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(8));
	CUT_6359:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(9));
	CUT_6360:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(10));
	CUT_6361:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(11));
	CUT_6362:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(12));
	CUT_6363:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(13));
	CUT_6364:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(14));
	CUT_6365:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(15));
	CUT_6366:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(16));
	CUT_6367:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(17));
	CUT_6368:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(18));
	CUT_6369:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(19));
	CUT_6370:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(20));
	CUT_6371:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(21));
	CUT_6372:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(22));
	CUT_6373:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(23));
	CUT_6374:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(24));
	CUT_6375:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(25));
	CUT_6376:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(26));
	CUT_6377:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(27));
	CUT_6378:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(28));
	CUT_6379:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(29));
	CUT_6380:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(30));
	CUT_6381:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(31));
	CUT_6382:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(32));
	CUT_6383:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(33));
	CUT_6384:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(34));
	CUT_6385:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(35));
	CUT_6386:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(36));
	CUT_6387:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(37));
	CUT_6388:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(38));
	CUT_6389:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(39));
	CUT_6390:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(40));
	CUT_6391:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(41));
	CUT_6392:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(42));
	CUT_6393:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(43));
	CUT_6394:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(44));
	CUT_6395:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(45));
	CUT_6396:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(46));
	CUT_6397:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(47));
	CUT_6398:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(48));
	CUT_6399:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(127)(49));
	CUT_6400:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(0));
	CUT_6401:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(1));
	CUT_6402:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(2));
	CUT_6403:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(3));
	CUT_6404:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(4));
	CUT_6405:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(5));
	CUT_6406:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(6));
	CUT_6407:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(7));
	CUT_6408:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(8));
	CUT_6409:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(9));
	CUT_6410:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(10));
	CUT_6411:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(11));
	CUT_6412:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(12));
	CUT_6413:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(13));
	CUT_6414:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(14));
	CUT_6415:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(15));
	CUT_6416:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(16));
	CUT_6417:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(17));
	CUT_6418:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(18));
	CUT_6419:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(19));
	CUT_6420:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(20));
	CUT_6421:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(21));
	CUT_6422:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(22));
	CUT_6423:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(23));
	CUT_6424:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(24));
	CUT_6425:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(25));
	CUT_6426:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(26));
	CUT_6427:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(27));
	CUT_6428:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(28));
	CUT_6429:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(29));
	CUT_6430:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(30));
	CUT_6431:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(31));
	CUT_6432:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(32));
	CUT_6433:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(33));
	CUT_6434:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(34));
	CUT_6435:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(35));
	CUT_6436:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(36));
	CUT_6437:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(37));
	CUT_6438:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(38));
	CUT_6439:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(39));
	CUT_6440:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(40));
	CUT_6441:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(41));
	CUT_6442:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(42));
	CUT_6443:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(43));
	CUT_6444:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(44));
	CUT_6445:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(45));
	CUT_6446:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(46));
	CUT_6447:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(47));
	CUT_6448:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(48));
	CUT_6449:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(128)(49));
	CUT_6450:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(0));
	CUT_6451:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(1));
	CUT_6452:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(2));
	CUT_6453:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(3));
	CUT_6454:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(4));
	CUT_6455:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(5));
	CUT_6456:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(6));
	CUT_6457:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(7));
	CUT_6458:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(8));
	CUT_6459:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(9));
	CUT_6460:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(10));
	CUT_6461:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(11));
	CUT_6462:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(12));
	CUT_6463:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(13));
	CUT_6464:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(14));
	CUT_6465:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(15));
	CUT_6466:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(16));
	CUT_6467:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(17));
	CUT_6468:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(18));
	CUT_6469:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(19));
	CUT_6470:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(20));
	CUT_6471:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(21));
	CUT_6472:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(22));
	CUT_6473:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(23));
	CUT_6474:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(24));
	CUT_6475:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(25));
	CUT_6476:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(26));
	CUT_6477:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(27));
	CUT_6478:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(28));
	CUT_6479:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(29));
	CUT_6480:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(30));
	CUT_6481:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(31));
	CUT_6482:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(32));
	CUT_6483:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(33));
	CUT_6484:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(34));
	CUT_6485:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(35));
	CUT_6486:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(36));
	CUT_6487:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(37));
	CUT_6488:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(38));
	CUT_6489:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(39));
	CUT_6490:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(40));
	CUT_6491:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(41));
	CUT_6492:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(42));
	CUT_6493:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(43));
	CUT_6494:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(44));
	CUT_6495:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(45));
	CUT_6496:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(46));
	CUT_6497:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(47));
	CUT_6498:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(48));
	CUT_6499:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(129)(49));
	CUT_6500:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(0));
	CUT_6501:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(1));
	CUT_6502:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(2));
	CUT_6503:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(3));
	CUT_6504:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(4));
	CUT_6505:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(5));
	CUT_6506:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(6));
	CUT_6507:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(7));
	CUT_6508:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(8));
	CUT_6509:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(9));
	CUT_6510:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(10));
	CUT_6511:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(11));
	CUT_6512:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(12));
	CUT_6513:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(13));
	CUT_6514:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(14));
	CUT_6515:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(15));
	CUT_6516:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(16));
	CUT_6517:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(17));
	CUT_6518:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(18));
	CUT_6519:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(19));
	CUT_6520:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(20));
	CUT_6521:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(21));
	CUT_6522:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(22));
	CUT_6523:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(23));
	CUT_6524:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(24));
	CUT_6525:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(25));
	CUT_6526:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(26));
	CUT_6527:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(27));
	CUT_6528:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(28));
	CUT_6529:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(29));
	CUT_6530:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(30));
	CUT_6531:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(31));
	CUT_6532:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(32));
	CUT_6533:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(33));
	CUT_6534:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(34));
	CUT_6535:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(35));
	CUT_6536:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(36));
	CUT_6537:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(37));
	CUT_6538:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(38));
	CUT_6539:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(39));
	CUT_6540:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(40));
	CUT_6541:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(41));
	CUT_6542:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(42));
	CUT_6543:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(43));
	CUT_6544:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(44));
	CUT_6545:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(45));
	CUT_6546:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(46));
	CUT_6547:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(47));
	CUT_6548:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(48));
	CUT_6549:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(130)(49));
	CUT_6550:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(0));
	CUT_6551:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(1));
	CUT_6552:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(2));
	CUT_6553:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(3));
	CUT_6554:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(4));
	CUT_6555:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(5));
	CUT_6556:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(6));
	CUT_6557:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(7));
	CUT_6558:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(8));
	CUT_6559:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(9));
	CUT_6560:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(10));
	CUT_6561:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(11));
	CUT_6562:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(12));
	CUT_6563:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(13));
	CUT_6564:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(14));
	CUT_6565:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(15));
	CUT_6566:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(16));
	CUT_6567:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(17));
	CUT_6568:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(18));
	CUT_6569:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(19));
	CUT_6570:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(20));
	CUT_6571:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(21));
	CUT_6572:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(22));
	CUT_6573:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(23));
	CUT_6574:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(24));
	CUT_6575:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(25));
	CUT_6576:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(26));
	CUT_6577:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(27));
	CUT_6578:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(28));
	CUT_6579:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(29));
	CUT_6580:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(30));
	CUT_6581:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(31));
	CUT_6582:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(32));
	CUT_6583:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(33));
	CUT_6584:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(34));
	CUT_6585:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(35));
	CUT_6586:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(36));
	CUT_6587:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(37));
	CUT_6588:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(38));
	CUT_6589:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(39));
	CUT_6590:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(40));
	CUT_6591:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(41));
	CUT_6592:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(42));
	CUT_6593:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(43));
	CUT_6594:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(44));
	CUT_6595:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(45));
	CUT_6596:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(46));
	CUT_6597:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(47));
	CUT_6598:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(48));
	CUT_6599:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(131)(49));
	CUT_6600:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(0));
	CUT_6601:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(1));
	CUT_6602:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(2));
	CUT_6603:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(3));
	CUT_6604:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(4));
	CUT_6605:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(5));
	CUT_6606:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(6));
	CUT_6607:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(7));
	CUT_6608:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(8));
	CUT_6609:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(9));
	CUT_6610:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(10));
	CUT_6611:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(11));
	CUT_6612:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(12));
	CUT_6613:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(13));
	CUT_6614:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(14));
	CUT_6615:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(15));
	CUT_6616:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(16));
	CUT_6617:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(17));
	CUT_6618:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(18));
	CUT_6619:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(19));
	CUT_6620:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(20));
	CUT_6621:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(21));
	CUT_6622:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(22));
	CUT_6623:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(23));
	CUT_6624:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(24));
	CUT_6625:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(25));
	CUT_6626:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(26));
	CUT_6627:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(27));
	CUT_6628:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(28));
	CUT_6629:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(29));
	CUT_6630:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(30));
	CUT_6631:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(31));
	CUT_6632:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(32));
	CUT_6633:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(33));
	CUT_6634:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(34));
	CUT_6635:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(35));
	CUT_6636:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(36));
	CUT_6637:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(37));
	CUT_6638:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(38));
	CUT_6639:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(39));
	CUT_6640:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(40));
	CUT_6641:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(41));
	CUT_6642:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(42));
	CUT_6643:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(43));
	CUT_6644:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(44));
	CUT_6645:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(45));
	CUT_6646:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(46));
	CUT_6647:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(47));
	CUT_6648:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(48));
	CUT_6649:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(132)(49));
	CUT_6650:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(0));
	CUT_6651:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(1));
	CUT_6652:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(2));
	CUT_6653:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(3));
	CUT_6654:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(4));
	CUT_6655:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(5));
	CUT_6656:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(6));
	CUT_6657:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(7));
	CUT_6658:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(8));
	CUT_6659:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(9));
	CUT_6660:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(10));
	CUT_6661:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(11));
	CUT_6662:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(12));
	CUT_6663:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(13));
	CUT_6664:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(14));
	CUT_6665:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(15));
	CUT_6666:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(16));
	CUT_6667:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(17));
	CUT_6668:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(18));
	CUT_6669:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(19));
	CUT_6670:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(20));
	CUT_6671:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(21));
	CUT_6672:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(22));
	CUT_6673:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(23));
	CUT_6674:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(24));
	CUT_6675:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(25));
	CUT_6676:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(26));
	CUT_6677:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(27));
	CUT_6678:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(28));
	CUT_6679:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(29));
	CUT_6680:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(30));
	CUT_6681:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(31));
	CUT_6682:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(32));
	CUT_6683:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(33));
	CUT_6684:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(34));
	CUT_6685:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(35));
	CUT_6686:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(36));
	CUT_6687:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(37));
	CUT_6688:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(38));
	CUT_6689:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(39));
	CUT_6690:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(40));
	CUT_6691:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(41));
	CUT_6692:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(42));
	CUT_6693:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(43));
	CUT_6694:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(44));
	CUT_6695:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(45));
	CUT_6696:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(46));
	CUT_6697:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(47));
	CUT_6698:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(48));
	CUT_6699:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(133)(49));
	CUT_6700:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(0));
	CUT_6701:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(1));
	CUT_6702:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(2));
	CUT_6703:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(3));
	CUT_6704:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(4));
	CUT_6705:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(5));
	CUT_6706:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(6));
	CUT_6707:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(7));
	CUT_6708:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(8));
	CUT_6709:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(9));
	CUT_6710:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(10));
	CUT_6711:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(11));
	CUT_6712:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(12));
	CUT_6713:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(13));
	CUT_6714:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(14));
	CUT_6715:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(15));
	CUT_6716:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(16));
	CUT_6717:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(17));
	CUT_6718:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(18));
	CUT_6719:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(19));
	CUT_6720:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(20));
	CUT_6721:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(21));
	CUT_6722:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(22));
	CUT_6723:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(23));
	CUT_6724:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(24));
	CUT_6725:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(25));
	CUT_6726:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(26));
	CUT_6727:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(27));
	CUT_6728:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(28));
	CUT_6729:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(29));
	CUT_6730:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(30));
	CUT_6731:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(31));
	CUT_6732:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(32));
	CUT_6733:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(33));
	CUT_6734:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(34));
	CUT_6735:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(35));
	CUT_6736:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(36));
	CUT_6737:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(37));
	CUT_6738:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(38));
	CUT_6739:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(39));
	CUT_6740:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(40));
	CUT_6741:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(41));
	CUT_6742:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(42));
	CUT_6743:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(43));
	CUT_6744:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(44));
	CUT_6745:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(45));
	CUT_6746:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(46));
	CUT_6747:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(47));
	CUT_6748:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(48));
	CUT_6749:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(134)(49));
	CUT_6750:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(0));
	CUT_6751:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(1));
	CUT_6752:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(2));
	CUT_6753:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(3));
	CUT_6754:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(4));
	CUT_6755:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(5));
	CUT_6756:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(6));
	CUT_6757:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(7));
	CUT_6758:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(8));
	CUT_6759:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(9));
	CUT_6760:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(10));
	CUT_6761:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(11));
	CUT_6762:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(12));
	CUT_6763:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(13));
	CUT_6764:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(14));
	CUT_6765:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(15));
	CUT_6766:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(16));
	CUT_6767:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(17));
	CUT_6768:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(18));
	CUT_6769:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(19));
	CUT_6770:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(20));
	CUT_6771:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(21));
	CUT_6772:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(22));
	CUT_6773:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(23));
	CUT_6774:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(24));
	CUT_6775:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(25));
	CUT_6776:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(26));
	CUT_6777:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(27));
	CUT_6778:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(28));
	CUT_6779:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(29));
	CUT_6780:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(30));
	CUT_6781:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(31));
	CUT_6782:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(32));
	CUT_6783:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(33));
	CUT_6784:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(34));
	CUT_6785:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(35));
	CUT_6786:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(36));
	CUT_6787:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(37));
	CUT_6788:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(38));
	CUT_6789:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(39));
	CUT_6790:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(40));
	CUT_6791:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(41));
	CUT_6792:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(42));
	CUT_6793:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(43));
	CUT_6794:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(44));
	CUT_6795:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(45));
	CUT_6796:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(46));
	CUT_6797:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(47));
	CUT_6798:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(48));
	CUT_6799:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(135)(49));
	CUT_6800:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(0));
	CUT_6801:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(1));
	CUT_6802:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(2));
	CUT_6803:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(3));
	CUT_6804:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(4));
	CUT_6805:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(5));
	CUT_6806:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(6));
	CUT_6807:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(7));
	CUT_6808:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(8));
	CUT_6809:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(9));
	CUT_6810:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(10));
	CUT_6811:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(11));
	CUT_6812:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(12));
	CUT_6813:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(13));
	CUT_6814:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(14));
	CUT_6815:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(15));
	CUT_6816:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(16));
	CUT_6817:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(17));
	CUT_6818:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(18));
	CUT_6819:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(19));
	CUT_6820:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(20));
	CUT_6821:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(21));
	CUT_6822:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(22));
	CUT_6823:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(23));
	CUT_6824:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(24));
	CUT_6825:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(25));
	CUT_6826:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(26));
	CUT_6827:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(27));
	CUT_6828:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(28));
	CUT_6829:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(29));
	CUT_6830:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(30));
	CUT_6831:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(31));
	CUT_6832:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(32));
	CUT_6833:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(33));
	CUT_6834:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(34));
	CUT_6835:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(35));
	CUT_6836:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(36));
	CUT_6837:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(37));
	CUT_6838:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(38));
	CUT_6839:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(39));
	CUT_6840:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(40));
	CUT_6841:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(41));
	CUT_6842:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(42));
	CUT_6843:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(43));
	CUT_6844:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(44));
	CUT_6845:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(45));
	CUT_6846:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(46));
	CUT_6847:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(47));
	CUT_6848:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(48));
	CUT_6849:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(136)(49));
	CUT_6850:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(0));
	CUT_6851:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(1));
	CUT_6852:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(2));
	CUT_6853:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(3));
	CUT_6854:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(4));
	CUT_6855:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(5));
	CUT_6856:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(6));
	CUT_6857:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(7));
	CUT_6858:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(8));
	CUT_6859:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(9));
	CUT_6860:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(10));
	CUT_6861:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(11));
	CUT_6862:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(12));
	CUT_6863:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(13));
	CUT_6864:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(14));
	CUT_6865:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(15));
	CUT_6866:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(16));
	CUT_6867:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(17));
	CUT_6868:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(18));
	CUT_6869:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(19));
	CUT_6870:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(20));
	CUT_6871:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(21));
	CUT_6872:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(22));
	CUT_6873:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(23));
	CUT_6874:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(24));
	CUT_6875:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(25));
	CUT_6876:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(26));
	CUT_6877:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(27));
	CUT_6878:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(28));
	CUT_6879:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(29));
	CUT_6880:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(30));
	CUT_6881:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(31));
	CUT_6882:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(32));
	CUT_6883:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(33));
	CUT_6884:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(34));
	CUT_6885:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(35));
	CUT_6886:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(36));
	CUT_6887:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(37));
	CUT_6888:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(38));
	CUT_6889:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(39));
	CUT_6890:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(40));
	CUT_6891:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(41));
	CUT_6892:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(42));
	CUT_6893:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(43));
	CUT_6894:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(44));
	CUT_6895:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(45));
	CUT_6896:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(46));
	CUT_6897:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(47));
	CUT_6898:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(48));
	CUT_6899:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(137)(49));
	CUT_6900:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(0));
	CUT_6901:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(1));
	CUT_6902:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(2));
	CUT_6903:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(3));
	CUT_6904:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(4));
	CUT_6905:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(5));
	CUT_6906:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(6));
	CUT_6907:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(7));
	CUT_6908:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(8));
	CUT_6909:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(9));
	CUT_6910:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(10));
	CUT_6911:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(11));
	CUT_6912:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(12));
	CUT_6913:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(13));
	CUT_6914:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(14));
	CUT_6915:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(15));
	CUT_6916:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(16));
	CUT_6917:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(17));
	CUT_6918:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(18));
	CUT_6919:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(19));
	CUT_6920:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(20));
	CUT_6921:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(21));
	CUT_6922:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(22));
	CUT_6923:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(23));
	CUT_6924:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(24));
	CUT_6925:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(25));
	CUT_6926:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(26));
	CUT_6927:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(27));
	CUT_6928:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(28));
	CUT_6929:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(29));
	CUT_6930:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(30));
	CUT_6931:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(31));
	CUT_6932:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(32));
	CUT_6933:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(33));
	CUT_6934:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(34));
	CUT_6935:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(35));
	CUT_6936:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(36));
	CUT_6937:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(37));
	CUT_6938:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(38));
	CUT_6939:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(39));
	CUT_6940:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(40));
	CUT_6941:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(41));
	CUT_6942:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(42));
	CUT_6943:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(43));
	CUT_6944:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(44));
	CUT_6945:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(45));
	CUT_6946:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(46));
	CUT_6947:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(47));
	CUT_6948:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(48));
	CUT_6949:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(138)(49));
	CUT_6950:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(0));
	CUT_6951:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(1));
	CUT_6952:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(2));
	CUT_6953:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(3));
	CUT_6954:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(4));
	CUT_6955:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(5));
	CUT_6956:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(6));
	CUT_6957:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(7));
	CUT_6958:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(8));
	CUT_6959:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(9));
	CUT_6960:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(10));
	CUT_6961:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(11));
	CUT_6962:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(12));
	CUT_6963:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(13));
	CUT_6964:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(14));
	CUT_6965:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(15));
	CUT_6966:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(16));
	CUT_6967:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(17));
	CUT_6968:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(18));
	CUT_6969:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(19));
	CUT_6970:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(20));
	CUT_6971:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(21));
	CUT_6972:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(22));
	CUT_6973:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(23));
	CUT_6974:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(24));
	CUT_6975:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(25));
	CUT_6976:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(26));
	CUT_6977:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(27));
	CUT_6978:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(28));
	CUT_6979:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(29));
	CUT_6980:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(30));
	CUT_6981:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(31));
	CUT_6982:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(32));
	CUT_6983:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(33));
	CUT_6984:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(34));
	CUT_6985:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(35));
	CUT_6986:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(36));
	CUT_6987:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(37));
	CUT_6988:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(38));
	CUT_6989:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(39));
	CUT_6990:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(40));
	CUT_6991:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(41));
	CUT_6992:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(42));
	CUT_6993:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(43));
	CUT_6994:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(44));
	CUT_6995:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(45));
	CUT_6996:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(46));
	CUT_6997:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(47));
	CUT_6998:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(48));
	CUT_6999:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(139)(49));
	CUT_7000:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(0));
	CUT_7001:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(1));
	CUT_7002:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(2));
	CUT_7003:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(3));
	CUT_7004:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(4));
	CUT_7005:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(5));
	CUT_7006:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(6));
	CUT_7007:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(7));
	CUT_7008:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(8));
	CUT_7009:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(9));
	CUT_7010:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(10));
	CUT_7011:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(11));
	CUT_7012:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(12));
	CUT_7013:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(13));
	CUT_7014:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(14));
	CUT_7015:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(15));
	CUT_7016:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(16));
	CUT_7017:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(17));
	CUT_7018:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(18));
	CUT_7019:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(19));
	CUT_7020:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(20));
	CUT_7021:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(21));
	CUT_7022:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(22));
	CUT_7023:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(23));
	CUT_7024:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(24));
	CUT_7025:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(25));
	CUT_7026:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(26));
	CUT_7027:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(27));
	CUT_7028:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(28));
	CUT_7029:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(29));
	CUT_7030:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(30));
	CUT_7031:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(31));
	CUT_7032:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(32));
	CUT_7033:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(33));
	CUT_7034:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(34));
	CUT_7035:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(35));
	CUT_7036:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(36));
	CUT_7037:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(37));
	CUT_7038:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(38));
	CUT_7039:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(39));
	CUT_7040:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(40));
	CUT_7041:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(41));
	CUT_7042:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(42));
	CUT_7043:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(43));
	CUT_7044:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(44));
	CUT_7045:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(45));
	CUT_7046:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(46));
	CUT_7047:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(47));
	CUT_7048:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(48));
	CUT_7049:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(140)(49));
	CUT_7050:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(0));
	CUT_7051:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(1));
	CUT_7052:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(2));
	CUT_7053:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(3));
	CUT_7054:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(4));
	CUT_7055:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(5));
	CUT_7056:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(6));
	CUT_7057:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(7));
	CUT_7058:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(8));
	CUT_7059:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(9));
	CUT_7060:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(10));
	CUT_7061:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(11));
	CUT_7062:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(12));
	CUT_7063:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(13));
	CUT_7064:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(14));
	CUT_7065:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(15));
	CUT_7066:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(16));
	CUT_7067:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(17));
	CUT_7068:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(18));
	CUT_7069:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(19));
	CUT_7070:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(20));
	CUT_7071:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(21));
	CUT_7072:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(22));
	CUT_7073:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(23));
	CUT_7074:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(24));
	CUT_7075:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(25));
	CUT_7076:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(26));
	CUT_7077:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(27));
	CUT_7078:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(28));
	CUT_7079:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(29));
	CUT_7080:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(30));
	CUT_7081:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(31));
	CUT_7082:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(32));
	CUT_7083:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(33));
	CUT_7084:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(34));
	CUT_7085:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(35));
	CUT_7086:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(36));
	CUT_7087:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(37));
	CUT_7088:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(38));
	CUT_7089:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(39));
	CUT_7090:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(40));
	CUT_7091:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(41));
	CUT_7092:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(42));
	CUT_7093:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(43));
	CUT_7094:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(44));
	CUT_7095:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(45));
	CUT_7096:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(46));
	CUT_7097:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(47));
	CUT_7098:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(48));
	CUT_7099:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(141)(49));
	CUT_7100:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(0));
	CUT_7101:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(1));
	CUT_7102:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(2));
	CUT_7103:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(3));
	CUT_7104:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(4));
	CUT_7105:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(5));
	CUT_7106:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(6));
	CUT_7107:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(7));
	CUT_7108:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(8));
	CUT_7109:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(9));
	CUT_7110:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(10));
	CUT_7111:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(11));
	CUT_7112:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(12));
	CUT_7113:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(13));
	CUT_7114:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(14));
	CUT_7115:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(15));
	CUT_7116:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(16));
	CUT_7117:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(17));
	CUT_7118:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(18));
	CUT_7119:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(19));
	CUT_7120:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(20));
	CUT_7121:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(21));
	CUT_7122:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(22));
	CUT_7123:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(23));
	CUT_7124:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(24));
	CUT_7125:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(25));
	CUT_7126:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(26));
	CUT_7127:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(27));
	CUT_7128:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(28));
	CUT_7129:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(29));
	CUT_7130:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(30));
	CUT_7131:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(31));
	CUT_7132:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(32));
	CUT_7133:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(33));
	CUT_7134:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(34));
	CUT_7135:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(35));
	CUT_7136:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(36));
	CUT_7137:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(37));
	CUT_7138:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(38));
	CUT_7139:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(39));
	CUT_7140:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(40));
	CUT_7141:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(41));
	CUT_7142:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(42));
	CUT_7143:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(43));
	CUT_7144:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(44));
	CUT_7145:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(45));
	CUT_7146:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(46));
	CUT_7147:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(47));
	CUT_7148:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(48));
	CUT_7149:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(142)(49));
	CUT_7150:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(0));
	CUT_7151:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(1));
	CUT_7152:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(2));
	CUT_7153:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(3));
	CUT_7154:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(4));
	CUT_7155:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(5));
	CUT_7156:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(6));
	CUT_7157:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(7));
	CUT_7158:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(8));
	CUT_7159:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(9));
	CUT_7160:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(10));
	CUT_7161:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(11));
	CUT_7162:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(12));
	CUT_7163:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(13));
	CUT_7164:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(14));
	CUT_7165:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(15));
	CUT_7166:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(16));
	CUT_7167:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(17));
	CUT_7168:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(18));
	CUT_7169:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(19));
	CUT_7170:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(20));
	CUT_7171:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(21));
	CUT_7172:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(22));
	CUT_7173:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(23));
	CUT_7174:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(24));
	CUT_7175:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(25));
	CUT_7176:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(26));
	CUT_7177:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(27));
	CUT_7178:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(28));
	CUT_7179:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(29));
	CUT_7180:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(30));
	CUT_7181:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(31));
	CUT_7182:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(32));
	CUT_7183:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(33));
	CUT_7184:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(34));
	CUT_7185:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(35));
	CUT_7186:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(36));
	CUT_7187:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(37));
	CUT_7188:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(38));
	CUT_7189:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(39));
	CUT_7190:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(40));
	CUT_7191:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(41));
	CUT_7192:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(42));
	CUT_7193:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(43));
	CUT_7194:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(44));
	CUT_7195:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(45));
	CUT_7196:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(46));
	CUT_7197:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(47));
	CUT_7198:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(48));
	CUT_7199:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(143)(49));
	CUT_7200:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(0));
	CUT_7201:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(1));
	CUT_7202:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(2));
	CUT_7203:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(3));
	CUT_7204:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(4));
	CUT_7205:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(5));
	CUT_7206:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(6));
	CUT_7207:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(7));
	CUT_7208:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(8));
	CUT_7209:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(9));
	CUT_7210:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(10));
	CUT_7211:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(11));
	CUT_7212:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(12));
	CUT_7213:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(13));
	CUT_7214:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(14));
	CUT_7215:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(15));
	CUT_7216:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(16));
	CUT_7217:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(17));
	CUT_7218:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(18));
	CUT_7219:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(19));
	CUT_7220:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(20));
	CUT_7221:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(21));
	CUT_7222:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(22));
	CUT_7223:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(23));
	CUT_7224:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(24));
	CUT_7225:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(25));
	CUT_7226:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(26));
	CUT_7227:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(27));
	CUT_7228:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(28));
	CUT_7229:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(29));
	CUT_7230:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(30));
	CUT_7231:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(31));
	CUT_7232:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(32));
	CUT_7233:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(33));
	CUT_7234:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(34));
	CUT_7235:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(35));
	CUT_7236:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(36));
	CUT_7237:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(37));
	CUT_7238:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(38));
	CUT_7239:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(39));
	CUT_7240:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(40));
	CUT_7241:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(41));
	CUT_7242:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(42));
	CUT_7243:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(43));
	CUT_7244:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(44));
	CUT_7245:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(45));
	CUT_7246:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(46));
	CUT_7247:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(47));
	CUT_7248:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(48));
	CUT_7249:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(144)(49));
	CUT_7250:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(0));
	CUT_7251:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(1));
	CUT_7252:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(2));
	CUT_7253:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(3));
	CUT_7254:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(4));
	CUT_7255:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(5));
	CUT_7256:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(6));
	CUT_7257:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(7));
	CUT_7258:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(8));
	CUT_7259:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(9));
	CUT_7260:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(10));
	CUT_7261:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(11));
	CUT_7262:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(12));
	CUT_7263:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(13));
	CUT_7264:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(14));
	CUT_7265:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(15));
	CUT_7266:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(16));
	CUT_7267:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(17));
	CUT_7268:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(18));
	CUT_7269:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(19));
	CUT_7270:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(20));
	CUT_7271:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(21));
	CUT_7272:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(22));
	CUT_7273:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(23));
	CUT_7274:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(24));
	CUT_7275:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(25));
	CUT_7276:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(26));
	CUT_7277:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(27));
	CUT_7278:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(28));
	CUT_7279:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(29));
	CUT_7280:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(30));
	CUT_7281:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(31));
	CUT_7282:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(32));
	CUT_7283:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(33));
	CUT_7284:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(34));
	CUT_7285:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(35));
	CUT_7286:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(36));
	CUT_7287:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(37));
	CUT_7288:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(38));
	CUT_7289:	entity work.CUT_Buff
	generic map(g_Buffer => "11")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(39));
	CUT_7290:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(40));
	CUT_7291:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(41));
	CUT_7292:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(42));
	CUT_7293:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(43));
	CUT_7294:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(44));
	CUT_7295:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(45));
	CUT_7296:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(46));
	CUT_7297:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(47));
	CUT_7298:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(48));
	CUT_7299:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(145)(49));
	CUT_7300:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(0));
	CUT_7301:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(1));
	CUT_7302:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(2));
	CUT_7303:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(3));
	CUT_7304:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(4));
	CUT_7305:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(5));
	CUT_7306:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(6));
	CUT_7307:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(7));
	CUT_7308:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(8));
	CUT_7309:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(9));
	CUT_7310:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(10));
	CUT_7311:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(11));
	CUT_7312:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(12));
	CUT_7313:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(13));
	CUT_7314:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(14));
	CUT_7315:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(15));
	CUT_7316:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(16));
	CUT_7317:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(17));
	CUT_7318:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(18));
	CUT_7319:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(19));
	CUT_7320:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(20));
	CUT_7321:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(21));
	CUT_7322:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(22));
	CUT_7323:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(23));
	CUT_7324:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(24));
	CUT_7325:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(25));
	CUT_7326:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(26));
	CUT_7327:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(27));
	CUT_7328:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(28));
	CUT_7329:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(29));
	CUT_7330:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(30));
	CUT_7331:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(31));
	CUT_7332:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(32));
	CUT_7333:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(33));
	CUT_7334:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(34));
	CUT_7335:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(35));
	CUT_7336:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(36));
	CUT_7337:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(37));
	CUT_7338:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(38));
	CUT_7339:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(39));
	CUT_7340:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(40));
	CUT_7341:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(41));
	CUT_7342:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(42));
	CUT_7343:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(43));
	CUT_7344:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(44));
	CUT_7345:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(45));
	CUT_7346:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(46));
	CUT_7347:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(47));
	CUT_7348:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(48));
	CUT_7349:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(146)(49));
	CUT_7350:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(0));
	CUT_7351:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(1));
	CUT_7352:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(2));
	CUT_7353:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(3));
	CUT_7354:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(4));
	CUT_7355:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(5));
	CUT_7356:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(6));
	CUT_7357:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(7));
	CUT_7358:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(8));
	CUT_7359:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(9));
	CUT_7360:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(10));
	CUT_7361:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(11));
	CUT_7362:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(12));
	CUT_7363:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(13));
	CUT_7364:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(14));
	CUT_7365:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(15));
	CUT_7366:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(16));
	CUT_7367:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(17));
	CUT_7368:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(18));
	CUT_7369:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(19));
	CUT_7370:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(20));
	CUT_7371:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(21));
	CUT_7372:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(22));
	CUT_7373:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(23));
	CUT_7374:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(24));
	CUT_7375:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(25));
	CUT_7376:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(26));
	CUT_7377:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(27));
	CUT_7378:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(28));
	CUT_7379:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(29));
	CUT_7380:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(30));
	CUT_7381:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(31));
	CUT_7382:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(32));
	CUT_7383:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(33));
	CUT_7384:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(34));
	CUT_7385:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(35));
	CUT_7386:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(36));
	CUT_7387:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(37));
	CUT_7388:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(38));
	CUT_7389:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(39));
	CUT_7390:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(40));
	CUT_7391:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(41));
	CUT_7392:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(42));
	CUT_7393:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(43));
	CUT_7394:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(44));
	CUT_7395:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(45));
	CUT_7396:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(46));
	CUT_7397:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(47));
	CUT_7398:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(48));
	CUT_7399:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(147)(49));
	CUT_7400:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(0));
	CUT_7401:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(1));
	CUT_7402:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(2));
	CUT_7403:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(3));
	CUT_7404:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(4));
	CUT_7405:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(5));
	CUT_7406:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(6));
	CUT_7407:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(7));
	CUT_7408:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(8));
	CUT_7409:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(9));
	CUT_7410:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(10));
	CUT_7411:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(11));
	CUT_7412:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(12));
	CUT_7413:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(13));
	CUT_7414:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(14));
	CUT_7415:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(15));
	CUT_7416:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(16));
	CUT_7417:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(17));
	CUT_7418:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(18));
	CUT_7419:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(19));
	CUT_7420:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(20));
	CUT_7421:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(21));
	CUT_7422:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(22));
	CUT_7423:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(23));
	CUT_7424:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(24));
	CUT_7425:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(25));
	CUT_7426:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(26));
	CUT_7427:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(27));
	CUT_7428:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(28));
	CUT_7429:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(29));
	CUT_7430:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(30));
	CUT_7431:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(31));
	CUT_7432:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(32));
	CUT_7433:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(33));
	CUT_7434:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(34));
	CUT_7435:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(35));
	CUT_7436:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(36));
	CUT_7437:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(37));
	CUT_7438:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(38));
	CUT_7439:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(39));
	CUT_7440:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(40));
	CUT_7441:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(41));
	CUT_7442:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(42));
	CUT_7443:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(43));
	CUT_7444:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(44));
	CUT_7445:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(45));
	CUT_7446:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(46));
	CUT_7447:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(47));
	CUT_7448:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(48));
	CUT_7449:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(148)(49));
	CUT_7450:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(0));
	CUT_7451:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(1));
	CUT_7452:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(2));
	CUT_7453:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(3));
	CUT_7454:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(4));
	CUT_7455:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(5));
	CUT_7456:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(6));
	CUT_7457:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(7));
	CUT_7458:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(8));
	CUT_7459:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(9));
	CUT_7460:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(10));
	CUT_7461:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(11));
	CUT_7462:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(12));
	CUT_7463:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(13));
	CUT_7464:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(14));
	CUT_7465:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(15));
	CUT_7466:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(16));
	CUT_7467:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(17));
	CUT_7468:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(18));
	CUT_7469:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(19));
	CUT_7470:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(20));
	CUT_7471:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(21));
	CUT_7472:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(22));
	CUT_7473:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(23));
	CUT_7474:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(24));
	CUT_7475:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(25));
	CUT_7476:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(26));
	CUT_7477:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(27));
	CUT_7478:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(28));
	CUT_7479:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(29));
	CUT_7480:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(30));
	CUT_7481:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(31));
	CUT_7482:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(32));
	CUT_7483:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(33));
	CUT_7484:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(34));
	CUT_7485:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(35));
	CUT_7486:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(36));
	CUT_7487:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(37));
	CUT_7488:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(38));
	CUT_7489:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(39));
	CUT_7490:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(40));
	CUT_7491:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(41));
	CUT_7492:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(42));
	CUT_7493:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(43));
	CUT_7494:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(44));
	CUT_7495:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(45));
	CUT_7496:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(46));
	CUT_7497:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(47));
	CUT_7498:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(48));
	CUT_7499:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(149)(49));
	CUT_7500:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(0));
	CUT_7501:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(1));
	CUT_7502:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(2));
	CUT_7503:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(3));
	CUT_7504:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(4));
	CUT_7505:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(5));
	CUT_7506:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(6));
	CUT_7507:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(7));
	CUT_7508:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(8));
	CUT_7509:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(9));
	CUT_7510:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(10));
	CUT_7511:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(11));
	CUT_7512:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(12));
	CUT_7513:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(13));
	CUT_7514:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(14));
	CUT_7515:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(15));
	CUT_7516:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(16));
	CUT_7517:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(17));
	CUT_7518:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(18));
	CUT_7519:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(19));
	CUT_7520:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(20));
	CUT_7521:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(21));
	CUT_7522:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(22));
	CUT_7523:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(23));
	CUT_7524:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(24));
	CUT_7525:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(25));
	CUT_7526:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(26));
	CUT_7527:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(27));
	CUT_7528:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(28));
	CUT_7529:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(29));
	CUT_7530:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(30));
	CUT_7531:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(31));
	CUT_7532:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(32));
	CUT_7533:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(33));
	CUT_7534:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(34));
	CUT_7535:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(35));
	CUT_7536:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(36));
	CUT_7537:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(37));
	CUT_7538:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(38));
	CUT_7539:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(39));
	CUT_7540:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(40));
	CUT_7541:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(41));
	CUT_7542:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(42));
	CUT_7543:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(43));
	CUT_7544:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(44));
	CUT_7545:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(45));
	CUT_7546:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(46));
	CUT_7547:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(47));
	CUT_7548:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(48));
	CUT_7549:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(150)(49));
	CUT_7550:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(0));
	CUT_7551:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(1));
	CUT_7552:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(2));
	CUT_7553:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(3));
	CUT_7554:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(4));
	CUT_7555:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(5));
	CUT_7556:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(6));
	CUT_7557:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(7));
	CUT_7558:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(8));
	CUT_7559:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(9));
	CUT_7560:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(10));
	CUT_7561:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(11));
	CUT_7562:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(12));
	CUT_7563:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(13));
	CUT_7564:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(14));
	CUT_7565:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(15));
	CUT_7566:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(16));
	CUT_7567:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(17));
	CUT_7568:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(18));
	CUT_7569:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(19));
	CUT_7570:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(20));
	CUT_7571:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(21));
	CUT_7572:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(22));
	CUT_7573:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(23));
	CUT_7574:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(24));
	CUT_7575:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(25));
	CUT_7576:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(26));
	CUT_7577:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(27));
	CUT_7578:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(28));
	CUT_7579:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(29));
	CUT_7580:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(30));
	CUT_7581:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(31));
	CUT_7582:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(32));
	CUT_7583:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(33));
	CUT_7584:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(34));
	CUT_7585:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(35));
	CUT_7586:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(36));
	CUT_7587:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(37));
	CUT_7588:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(38));
	CUT_7589:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(39));
	CUT_7590:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(40));
	CUT_7591:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(41));
	CUT_7592:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(42));
	CUT_7593:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(43));
	CUT_7594:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(44));
	CUT_7595:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(45));
	CUT_7596:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(46));
	CUT_7597:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(47));
	CUT_7598:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(48));
	CUT_7599:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(151)(49));
	CUT_7600:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(0));
	CUT_7601:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(1));
	CUT_7602:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(2));
	CUT_7603:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(3));
	CUT_7604:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(4));
	CUT_7605:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(5));
	CUT_7606:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(6));
	CUT_7607:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(7));
	CUT_7608:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(8));
	CUT_7609:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(9));
	CUT_7610:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(10));
	CUT_7611:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(11));
	CUT_7612:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(12));
	CUT_7613:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(13));
	CUT_7614:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(14));
	CUT_7615:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(15));
	CUT_7616:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(16));
	CUT_7617:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(17));
	CUT_7618:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(18));
	CUT_7619:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(19));
	CUT_7620:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(20));
	CUT_7621:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(21));
	CUT_7622:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(22));
	CUT_7623:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(23));
	CUT_7624:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(24));
	CUT_7625:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(25));
	CUT_7626:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(26));
	CUT_7627:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(27));
	CUT_7628:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(28));
	CUT_7629:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(29));
	CUT_7630:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(30));
	CUT_7631:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(31));
	CUT_7632:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(32));
	CUT_7633:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(33));
	CUT_7634:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(34));
	CUT_7635:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(35));
	CUT_7636:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(36));
	CUT_7637:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(37));
	CUT_7638:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(38));
	CUT_7639:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(39));
	CUT_7640:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(40));
	CUT_7641:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(41));
	CUT_7642:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(42));
	CUT_7643:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(43));
	CUT_7644:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(44));
	CUT_7645:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(45));
	CUT_7646:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(46));
	CUT_7647:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(47));
	CUT_7648:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(48));
	CUT_7649:	entity work.CUT_Buff
	generic map(g_Buffer => "10")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(152)(49));
	CUT_7650:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(0));
	CUT_7651:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(1));
	CUT_7652:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(2));
	CUT_7653:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(3));
	CUT_7654:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(4));
	CUT_7655:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(5));
	CUT_7656:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(6));
	CUT_7657:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(7));
	CUT_7658:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(8));
	CUT_7659:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(9));
	CUT_7660:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(10));
	CUT_7661:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(11));
	CUT_7662:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(12));
	CUT_7663:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(13));
	CUT_7664:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(14));
	CUT_7665:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(15));
	CUT_7666:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(16));
	CUT_7667:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(17));
	CUT_7668:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(18));
	CUT_7669:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(19));
	CUT_7670:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(20));
	CUT_7671:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(21));
	CUT_7672:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(22));
	CUT_7673:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(23));
	CUT_7674:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(24));
	CUT_7675:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(25));
	CUT_7676:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(26));
	CUT_7677:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(27));
	CUT_7678:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(28));
	CUT_7679:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(29));
	CUT_7680:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(30));
	CUT_7681:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(31));
	CUT_7682:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(32));
	CUT_7683:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(33));
	CUT_7684:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(34));
	CUT_7685:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(35));
	CUT_7686:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(36));
	CUT_7687:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(37));
	CUT_7688:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(38));
	CUT_7689:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(39));
	CUT_7690:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(40));
	CUT_7691:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(41));
	CUT_7692:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(42));
	CUT_7693:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(43));
	CUT_7694:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(44));
	CUT_7695:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(45));
	CUT_7696:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(46));
	CUT_7697:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(47));
	CUT_7698:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(48));
	CUT_7699:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(153)(49));
	CUT_7700:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(0));
	CUT_7701:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(1));
	CUT_7702:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(2));
	CUT_7703:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(3));
	CUT_7704:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(4));
	CUT_7705:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(5));
	CUT_7706:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(6));
	CUT_7707:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(7));
	CUT_7708:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(8));
	CUT_7709:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(9));
	CUT_7710:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(10));
	CUT_7711:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(11));
	CUT_7712:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(12));
	CUT_7713:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(13));
	CUT_7714:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(14));
	CUT_7715:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(15));
	CUT_7716:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(16));
	CUT_7717:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(17));
	CUT_7718:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(18));
	CUT_7719:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(19));
	CUT_7720:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(20));
	CUT_7721:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(21));
	CUT_7722:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(22));
	CUT_7723:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(23));
	CUT_7724:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(24));
	CUT_7725:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(25));
	CUT_7726:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(26));
	CUT_7727:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(27));
	CUT_7728:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(28));
	CUT_7729:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(29));
	CUT_7730:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(30));
	CUT_7731:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(31));
	CUT_7732:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(32));
	CUT_7733:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(33));
	CUT_7734:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(34));
	CUT_7735:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(35));
	CUT_7736:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(36));
	CUT_7737:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(37));
	CUT_7738:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(38));
	CUT_7739:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(39));
	CUT_7740:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(40));
	CUT_7741:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(41));
	CUT_7742:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(42));
	CUT_7743:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(43));
	CUT_7744:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(44));
	CUT_7745:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(45));
	CUT_7746:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(46));
	CUT_7747:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(47));
	CUT_7748:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(48));
	CUT_7749:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(154)(49));
	CUT_7750:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(0));
	CUT_7751:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(1));
	CUT_7752:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(2));
	CUT_7753:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(3));
	CUT_7754:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(4));
	CUT_7755:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(5));
	CUT_7756:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(6));
	CUT_7757:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(7));
	CUT_7758:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(8));
	CUT_7759:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(9));
	CUT_7760:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(10));
	CUT_7761:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(11));
	CUT_7762:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(12));
	CUT_7763:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(13));
	CUT_7764:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(14));
	CUT_7765:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(15));
	CUT_7766:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(16));
	CUT_7767:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(17));
	CUT_7768:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(18));
	CUT_7769:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(19));
	CUT_7770:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(20));
	CUT_7771:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(21));
	CUT_7772:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(22));
	CUT_7773:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(23));
	CUT_7774:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(24));
	CUT_7775:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(25));
	CUT_7776:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(26));
	CUT_7777:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(27));
	CUT_7778:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(28));
	CUT_7779:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(29));
	CUT_7780:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(30));
	CUT_7781:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(31));
	CUT_7782:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(32));
	CUT_7783:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(33));
	CUT_7784:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(34));
	CUT_7785:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(35));
	CUT_7786:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(36));
	CUT_7787:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(37));
	CUT_7788:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(38));
	CUT_7789:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(39));
	CUT_7790:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(40));
	CUT_7791:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(41));
	CUT_7792:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(42));
	CUT_7793:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(43));
	CUT_7794:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(44));
	CUT_7795:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(45));
	CUT_7796:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(46));
	CUT_7797:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(47));
	CUT_7798:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(48));
	CUT_7799:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(155)(49));
	CUT_7800:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(0));
	CUT_7801:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(1));
	CUT_7802:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(2));
	CUT_7803:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(3));
	CUT_7804:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(4));
	CUT_7805:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(5));
	CUT_7806:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(6));
	CUT_7807:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(7));
	CUT_7808:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(8));
	CUT_7809:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(9));
	CUT_7810:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(10));
	CUT_7811:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(11));
	CUT_7812:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(12));
	CUT_7813:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(13));
	CUT_7814:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(14));
	CUT_7815:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(15));
	CUT_7816:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(16));
	CUT_7817:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(17));
	CUT_7818:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(18));
	CUT_7819:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(19));
	CUT_7820:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(20));
	CUT_7821:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(21));
	CUT_7822:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(22));
	CUT_7823:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(23));
	CUT_7824:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(24));
	CUT_7825:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(25));
	CUT_7826:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(26));
	CUT_7827:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(27));
	CUT_7828:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(28));
	CUT_7829:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(29));
	CUT_7830:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(30));
	CUT_7831:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(31));
	CUT_7832:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(32));
	CUT_7833:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(33));
	CUT_7834:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(34));
	CUT_7835:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(35));
	CUT_7836:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(36));
	CUT_7837:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(37));
	CUT_7838:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(38));
	CUT_7839:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(39));
	CUT_7840:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(40));
	CUT_7841:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(41));
	CUT_7842:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(42));
	CUT_7843:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(43));
	CUT_7844:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(44));
	CUT_7845:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(45));
	CUT_7846:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(46));
	CUT_7847:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(47));
	CUT_7848:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(48));
	CUT_7849:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(156)(49));
	CUT_7850:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(0));
	CUT_7851:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(1));
	CUT_7852:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(2));
	CUT_7853:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(3));
	CUT_7854:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(4));
	CUT_7855:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(5));
	CUT_7856:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(6));
	CUT_7857:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(7));
	CUT_7858:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(8));
	CUT_7859:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(9));
	CUT_7860:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(10));
	CUT_7861:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(11));
	CUT_7862:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(12));
	CUT_7863:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(13));
	CUT_7864:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(14));
	CUT_7865:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(15));
	CUT_7866:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(16));
	CUT_7867:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(17));
	CUT_7868:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(18));
	CUT_7869:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(19));
	CUT_7870:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(20));
	CUT_7871:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(21));
	CUT_7872:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(22));
	CUT_7873:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(23));
	CUT_7874:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(24));
	CUT_7875:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(25));
	CUT_7876:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(26));
	CUT_7877:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(27));
	CUT_7878:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(28));
	CUT_7879:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(29));
	CUT_7880:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(30));
	CUT_7881:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(31));
	CUT_7882:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(32));
	CUT_7883:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(33));
	CUT_7884:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(34));
	CUT_7885:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(35));
	CUT_7886:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(36));
	CUT_7887:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(37));
	CUT_7888:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(38));
	CUT_7889:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(39));
	CUT_7890:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(40));
	CUT_7891:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(41));
	CUT_7892:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(42));
	CUT_7893:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(43));
	CUT_7894:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(44));
	CUT_7895:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(45));
	CUT_7896:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(46));
	CUT_7897:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(47));
	CUT_7898:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(48));
	CUT_7899:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(157)(49));
	CUT_7900:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(0));
	CUT_7901:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(1));
	CUT_7902:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(2));
	CUT_7903:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(3));
	CUT_7904:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(4));
	CUT_7905:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(5));
	CUT_7906:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(6));
	CUT_7907:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(7));
	CUT_7908:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(8));
	CUT_7909:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(9));
	CUT_7910:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(10));
	CUT_7911:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(11));
	CUT_7912:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(12));
	CUT_7913:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(13));
	CUT_7914:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(14));
	CUT_7915:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(15));
	CUT_7916:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(16));
	CUT_7917:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(17));
	CUT_7918:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(18));
	CUT_7919:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(19));
	CUT_7920:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(20));
	CUT_7921:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(21));
	CUT_7922:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(22));
	CUT_7923:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(23));
	CUT_7924:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(24));
	CUT_7925:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(25));
	CUT_7926:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(26));
	CUT_7927:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(27));
	CUT_7928:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(28));
	CUT_7929:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(29));
	CUT_7930:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(30));
	CUT_7931:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(31));
	CUT_7932:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(32));
	CUT_7933:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(33));
	CUT_7934:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(34));
	CUT_7935:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(35));
	CUT_7936:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(36));
	CUT_7937:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(37));
	CUT_7938:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(38));
	CUT_7939:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(39));
	CUT_7940:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(40));
	CUT_7941:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(41));
	CUT_7942:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(42));
	CUT_7943:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(43));
	CUT_7944:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(44));
	CUT_7945:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(45));
	CUT_7946:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(46));
	CUT_7947:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(47));
	CUT_7948:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(48));
	CUT_7949:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(158)(49));
	CUT_7950:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(0));
	CUT_7951:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(1));
	CUT_7952:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(2));
	CUT_7953:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(3));
	CUT_7954:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(4));
	CUT_7955:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(5));
	CUT_7956:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(6));
	CUT_7957:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(7));
	CUT_7958:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(8));
	CUT_7959:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(9));
	CUT_7960:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(10));
	CUT_7961:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(11));
	CUT_7962:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(12));
	CUT_7963:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(13));
	CUT_7964:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(14));
	CUT_7965:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(15));
	CUT_7966:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(16));
	CUT_7967:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(17));
	CUT_7968:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(18));
	CUT_7969:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(19));
	CUT_7970:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(20));
	CUT_7971:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(21));
	CUT_7972:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(22));
	CUT_7973:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(23));
	CUT_7974:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(24));
	CUT_7975:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(25));
	CUT_7976:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(26));
	CUT_7977:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(27));
	CUT_7978:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(28));
	CUT_7979:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(29));
	CUT_7980:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(30));
	CUT_7981:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(31));
	CUT_7982:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(32));
	CUT_7983:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(33));
	CUT_7984:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(34));
	CUT_7985:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(35));
	CUT_7986:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(36));
	CUT_7987:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(37));
	CUT_7988:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(38));
	CUT_7989:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(39));
	CUT_7990:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(40));
	CUT_7991:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(41));
	CUT_7992:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(42));
	CUT_7993:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(43));
	CUT_7994:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(44));
	CUT_7995:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(45));
	CUT_7996:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(46));
	CUT_7997:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(47));
	CUT_7998:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(48));
	CUT_7999:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(159)(49));
	CUT_8000:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(0));
	CUT_8001:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(1));
	CUT_8002:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(2));
	CUT_8003:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(3));
	CUT_8004:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(4));
	CUT_8005:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(5));
	CUT_8006:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(6));
	CUT_8007:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(7));
	CUT_8008:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(8));
	CUT_8009:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(9));
	CUT_8010:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(10));
	CUT_8011:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(11));
	CUT_8012:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(12));
	CUT_8013:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(13));
	CUT_8014:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(14));
	CUT_8015:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(15));
	CUT_8016:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(16));
	CUT_8017:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(17));
	CUT_8018:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(18));
	CUT_8019:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(19));
	CUT_8020:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(20));
	CUT_8021:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(21));
	CUT_8022:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(22));
	CUT_8023:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(23));
	CUT_8024:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(24));
	CUT_8025:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(25));
	CUT_8026:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(26));
	CUT_8027:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(27));
	CUT_8028:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(28));
	CUT_8029:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(29));
	CUT_8030:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(30));
	CUT_8031:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(31));
	CUT_8032:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(32));
	CUT_8033:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(33));
	CUT_8034:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(34));
	CUT_8035:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(35));
	CUT_8036:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(36));
	CUT_8037:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(37));
	CUT_8038:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(38));
	CUT_8039:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(39));
	CUT_8040:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(40));
	CUT_8041:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(41));
	CUT_8042:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(42));
	CUT_8043:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(43));
	CUT_8044:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(44));
	CUT_8045:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(45));
	CUT_8046:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(46));
	CUT_8047:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(47));
	CUT_8048:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(48));
	CUT_8049:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(160)(49));
	CUT_8050:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(0));
	CUT_8051:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(1));
	CUT_8052:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(2));
	CUT_8053:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(3));
	CUT_8054:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(4));
	CUT_8055:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(5));
	CUT_8056:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(6));
	CUT_8057:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(7));
	CUT_8058:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(8));
	CUT_8059:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(9));
	CUT_8060:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(10));
	CUT_8061:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(11));
	CUT_8062:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(12));
	CUT_8063:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(13));
	CUT_8064:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(14));
	CUT_8065:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(15));
	CUT_8066:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(16));
	CUT_8067:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(17));
	CUT_8068:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(18));
	CUT_8069:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(19));
	CUT_8070:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(20));
	CUT_8071:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(21));
	CUT_8072:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(22));
	CUT_8073:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(23));
	CUT_8074:	entity work.CUT_Buff
	generic map(g_Buffer => "00")
	port map(i_Clk_Launch, i_Clk_Sample, i_CE, i_CLR, w_Error(161)(24));

	o_Error	<=	w_Error;

end architecture;